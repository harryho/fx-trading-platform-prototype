20101227,144000,1.5412,1.5412,1.5411,1.5412
20101227,144100,1.5413,1.5413,1.5413,1.5413
20101227,144200,1.5409,1.5409,1.5409,1.5409
20101227,144300,1.5409,1.5409,1.5409,1.5409
20101227,144400,1.5407,1.5407,1.5407,1.5407
20101227,144500,1.5408,1.5408,1.5408,1.5408
20101227,144700,1.5407,1.5407,1.5407,1.5407
20101227,144900,1.5409,1.5409,1.5409,1.5409
20101227,145100,1.541,1.541,1.5408,1.5408
20101227,145200,1.5408,1.5408,1.5407,1.5407
20101227,145300,1.5406,1.5406,1.5404,1.5404
20101227,145400,1.5404,1.5406,1.5404,1.5404
20101227,145500,1.5405,1.5406,1.5405,1.5406
20101227,145600,1.5407,1.5407,1.5407,1.5407
20101227,145800,1.541,1.541,1.541,1.541
20101227,150000,1.5412,1.5412,1.5412,1.5412
20101227,150100,1.5412,1.5412,1.5412,1.5412
20101227,150200,1.541,1.541,1.541,1.541
20101227,150300,1.5412,1.5412,1.5412,1.5412
20101227,150400,1.541,1.541,1.541,1.541
20101227,150500,1.5408,1.5408,1.5408,1.5408
20101227,150700,1.5409,1.5409,1.5409,1.5409
20101227,150900,1.5408,1.541,1.5408,1.541
20101227,151000,1.541,1.5411,1.541,1.541
20101227,151100,1.541,1.541,1.541,1.541
20101227,151300,1.5414,1.5414,1.5414,1.5414
20101227,151500,1.541,1.541,1.541,1.541
20101227,151700,1.5414,1.5414,1.5414,1.5414
20101227,151900,1.5414,1.5414,1.5414,1.5414
20101227,152000,1.5414,1.5414,1.5414,1.5414
20101227,152200,1.5413,1.5413,1.5413,1.5413
20101227,152400,1.5414,1.5414,1.5414,1.5414
20101227,152500,1.5414,1.5414,1.5414,1.5414
20101227,152700,1.5415,1.5415,1.5414,1.5415
20101227,152800,1.5413,1.5413,1.5413,1.5413
20101227,152900,1.5413,1.5413,1.5413,1.5413
20101227,153100,1.5412,1.5413,1.5412,1.5413
20101227,153200,1.5414,1.5415,1.5414,1.5414
20101227,153300,1.5413,1.5413,1.5413,1.5413
20101227,153500,1.5413,1.5413,1.5413,1.5413
20101227,153700,1.5409,1.5409,1.5409,1.5409
20101227,153900,1.5408,1.5408,1.5402,1.5402
20101227,154000,1.5403,1.5406,1.5403,1.5404
20101227,154100,1.5404,1.5405,1.5404,1.5404
20101227,154200,1.5404,1.5404,1.5404,1.5404
20101227,154400,1.5407,1.5407,1.5407,1.5407
20101227,154500,1.5408,1.5408,1.5408,1.5408
20101227,154600,1.5402,1.5402,1.5402,1.5402
20101227,154700,1.5402,1.5402,1.5402,1.5402
20101227,154800,1.5399,1.5399,1.5399,1.5399
20101227,155000,1.5401,1.5401,1.5401,1.5401
20101227,155200,1.5402,1.5403,1.5402,1.5403
20101227,155300,1.54,1.54,1.54,1.54
20101227,155400,1.5399,1.5399,1.5399,1.5399
20101227,155500,1.5397,1.5397,1.5397,1.5397
20101227,155600,1.5394,1.5394,1.5394,1.5394
20101227,155700,1.5394,1.5394,1.5394,1.5394
20101227,155900,1.5393,1.5393,1.5389,1.539
20101227,160000,1.5387,1.5387,1.5387,1.5387
20101227,160100,1.5388,1.5388,1.5388,1.5388
20101227,160300,1.539,1.539,1.539,1.539
20101227,160400,1.539,1.539,1.539,1.539
20101227,160500,1.5388,1.5388,1.5388,1.5388
20101227,160700,1.5389,1.5389,1.5387,1.5388
20101227,160800,1.5385,1.5385,1.5385,1.5385
20101227,161000,1.5384,1.5386,1.5384,1.5386
20101227,161100,1.5385,1.5387,1.5385,1.5387
20101227,161200,1.5387,1.5387,1.5387,1.5387
20101227,161400,1.5388,1.5388,1.5387,1.5387
20101227,161500,1.5386,1.5386,1.5383,1.5384
20101227,161600,1.5385,1.5385,1.5383,1.5384
20101227,161700,1.5383,1.5384,1.5383,1.5384
20101227,161800,1.5388,1.5388,1.5388,1.5388
20101227,162000,1.5384,1.5384,1.5384,1.5384
20101227,162100,1.5383,1.5383,1.5383,1.5383
20101227,162300,1.5382,1.5382,1.538,1.538
20101227,162400,1.5381,1.5381,1.5381,1.5381
20101227,162500,1.5381,1.5381,1.5381,1.5381
20101227,162600,1.538,1.538,1.538,1.538
20101227,162800,1.5378,1.5378,1.5378,1.5378
20101227,162900,1.5377,1.5377,1.5377,1.5377
20101227,163000,1.5373,1.5373,1.5373,1.5373
20101227,163100,1.5368,1.5368,1.5368,1.5368
20101227,163200,1.5369,1.5369,1.5369,1.5369
20101227,163300,1.5374,1.5374,1.5374,1.5374
20101227,163500,1.5377,1.5377,1.5377,1.5377
20101227,163600,1.5374,1.5374,1.5374,1.5374
20101227,163800,1.5373,1.5375,1.5373,1.5375
20101227,163900,1.5375,1.5375,1.5375,1.5375
20101227,164100,1.5372,1.5372,1.5372,1.5372
20101227,164200,1.5372,1.5372,1.5372,1.5372
20101227,164300,1.5372,1.5372,1.5372,1.5372
20101227,164500,1.5371,1.5373,1.5371,1.5373
20101227,164600,1.5375,1.5375,1.5375,1.5375
20101227,164700,1.5377,1.5377,1.5377,1.5377
20101227,164900,1.5375,1.5375,1.5375,1.5375
20101227,165100,1.5375,1.5375,1.5374,1.5374
20101227,165200,1.5375,1.5376,1.5375,1.5375
20101227,165300,1.5375,1.5375,1.5374,1.5375
20101227,165400,1.5377,1.5377,1.5377,1.5377
20101227,165500,1.5376,1.5376,1.5376,1.5376
20101227,165700,1.5377,1.5377,1.5377,1.5377
20101227,165900,1.5379,1.5379,1.5379,1.5379
20101227,170000,1.5379,1.5379,1.5379,1.5379
20101227,170200,1.5378,1.5378,1.5378,1.5378
20101227,170300,1.5378,1.5378,1.5378,1.5378
20101227,170400,1.5378,1.5378,1.5378,1.5378
20101227,170600,1.5378,1.5379,1.5378,1.5379
20101227,170700,1.538,1.538,1.538,1.538
20101227,170800,1.5381,1.5381,1.538,1.5381
20101227,170900,1.5381,1.5381,1.538,1.5381
20101227,171000,1.5381,1.5381,1.5381,1.5381
20101227,171200,1.5381,1.5381,1.5381,1.5381
20101227,171400,1.5381,1.5381,1.538,1.538
20101227,171500,1.5378,1.5378,1.5378,1.5378
20101227,171700,1.5378,1.5379,1.5378,1.5379
20101227,171800,1.5381,1.5381,1.5381,1.5381
20101227,171900,1.5381,1.5381,1.5381,1.5381
20101227,172100,1.5381,1.5381,1.5381,1.5381
20101227,172200,1.5381,1.5381,1.5381,1.5381
20101227,172300,1.5382,1.5382,1.5381,1.5381
20101227,172400,1.5382,1.5384,1.5382,1.5384
20101227,172500,1.5385,1.5385,1.5385,1.5385
20101227,172600,1.5385,1.5385,1.5385,1.5385
20101227,172800,1.5384,1.5384,1.5384,1.5384
20101227,173000,1.5385,1.5385,1.5385,1.5385
20101227,173100,1.5384,1.5384,1.5384,1.5384
20101227,173300,1.5385,1.5385,1.5383,1.5383
20101227,173400,1.5383,1.5383,1.5383,1.5383
20101227,173500,1.5385,1.5385,1.5385,1.5385
20101227,173600,1.5379,1.5379,1.5379,1.5379
20101227,173800,1.5379,1.5379,1.5379,1.5379
20101227,173900,1.538,1.5382,1.538,1.5381
20101227,174000,1.5381,1.5381,1.538,1.538
20101227,174100,1.5379,1.5381,1.5378,1.5381
20101227,174200,1.5381,1.5381,1.5381,1.5381
20101227,174300,1.538,1.538,1.538,1.538
20101227,174400,1.5379,1.5379,1.5379,1.5379
20101227,174500,1.5381,1.5381,1.5381,1.5381
20101227,174700,1.5381,1.5383,1.5381,1.5383
20101227,174800,1.5382,1.5382,1.5381,1.5382
20101227,174900,1.5381,1.5382,1.5381,1.5381
20101227,175000,1.5386,1.5386,1.5386,1.5386
20101227,175100,1.5385,1.5385,1.5385,1.5385
20101227,175200,1.5385,1.5385,1.5385,1.5385
20101227,175400,1.5385,1.5385,1.5385,1.5385
20101227,175500,1.5385,1.5386,1.5383,1.5386
20101227,175600,1.5386,1.5388,1.5386,1.5388
20101227,175700,1.5388,1.5392,1.5388,1.5392
20101227,175800,1.5393,1.5393,1.5393,1.5393
20101227,175900,1.5391,1.5391,1.5391,1.5391
20101227,180000,1.5392,1.5392,1.5388,1.5391
20101227,180100,1.5388,1.539,1.5386,1.5389
20101227,180200,1.539,1.539,1.5382,1.5383
20101227,180300,1.5382,1.5384,1.5382,1.5384
20101227,180400,1.5385,1.5389,1.5385,1.5389
20101227,180500,1.5389,1.5389,1.5387,1.5388
20101227,180600,1.5387,1.539,1.5387,1.5389
20101227,180700,1.5389,1.5391,1.5389,1.5391
20101227,180800,1.539,1.539,1.5389,1.539
20101227,180900,1.5389,1.5389,1.5388,1.5388
20101227,181000,1.5388,1.539,1.5388,1.539
20101227,181100,1.539,1.539,1.539,1.539
20101227,181200,1.539,1.5391,1.539,1.5391
20101227,181300,1.539,1.539,1.539,1.539
20101227,181400,1.5391,1.5394,1.539,1.5394
20101227,181500,1.5393,1.5394,1.5393,1.5393
20101227,181600,1.5393,1.5394,1.5393,1.5394
20101227,181700,1.5394,1.5395,1.5394,1.5395
20101227,181800,1.5395,1.5396,1.5395,1.5396
20101227,181900,1.5396,1.5396,1.5396,1.5396
20101227,182000,1.5396,1.5396,1.5396,1.5396
20101227,182100,1.5396,1.5398,1.5396,1.5398
20101227,182200,1.5399,1.5399,1.5399,1.5399
20101227,182300,1.5398,1.5398,1.5398,1.5398
20101227,182400,1.5398,1.5398,1.5397,1.5398
20101227,182500,1.5398,1.5398,1.5397,1.5398
20101227,182600,1.5398,1.5398,1.5397,1.5397
20101227,182700,1.5397,1.5399,1.5397,1.5399
20101227,182800,1.5399,1.5399,1.5398,1.5398
20101227,182900,1.5399,1.5399,1.5397,1.5397
20101227,183000,1.5398,1.5398,1.5396,1.5396
20101227,183100,1.5397,1.5397,1.5397,1.5397
20101227,183200,1.5397,1.5398,1.5397,1.5398
20101227,183300,1.5399,1.5399,1.5398,1.5398
20101227,183400,1.5398,1.5398,1.5397,1.5397
20101227,183500,1.5398,1.5398,1.5397,1.5397
20101227,183600,1.5397,1.5398,1.5397,1.5397
20101227,183700,1.5397,1.5397,1.5396,1.5397
20101227,183800,1.5397,1.5398,1.5396,1.5396
20101227,183900,1.5397,1.5397,1.5396,1.5396
20101227,184000,1.5396,1.5398,1.5396,1.5398
20101227,184100,1.5399,1.54,1.5399,1.54
20101227,184200,1.5399,1.54,1.5399,1.5399
20101227,184300,1.54,1.54,1.5398,1.5399
20101227,184400,1.5398,1.54,1.5398,1.5398
20101227,184500,1.5399,1.5404,1.5399,1.5404
20101227,184600,1.5403,1.5403,1.5401,1.5401
20101227,184700,1.5401,1.5401,1.5401,1.5401
20101227,184800,1.5402,1.5402,1.5402,1.5402
20101227,184900,1.5403,1.5403,1.5402,1.5403
20101227,185000,1.5404,1.5406,1.5404,1.5405
20101227,185100,1.5406,1.5406,1.5404,1.5404
20101227,185200,1.5405,1.5406,1.5404,1.5404
20101227,185300,1.5403,1.5403,1.5398,1.5398
20101227,185400,1.5399,1.54,1.5399,1.54
20101227,185500,1.5399,1.54,1.5399,1.54
20101227,185600,1.5401,1.5402,1.54,1.54
20101227,185700,1.54,1.54,1.5399,1.5399
20101227,185800,1.5399,1.54,1.5399,1.5399
20101227,185900,1.54,1.54,1.5399,1.5399
20101227,190000,1.5399,1.5399,1.5399,1.5399
20101227,190100,1.54,1.54,1.5398,1.5398
20101227,190200,1.5398,1.5398,1.5397,1.5398
20101227,190300,1.5398,1.5399,1.5398,1.5399
20101227,190400,1.5398,1.5398,1.5397,1.5397
20101227,190500,1.5398,1.5399,1.5398,1.5399
20101227,190600,1.5399,1.5399,1.5398,1.5399
20101227,190700,1.5399,1.5399,1.5397,1.5398
20101227,190800,1.5399,1.5401,1.5399,1.5401
20101227,190900,1.5401,1.5401,1.5401,1.5401
20101227,191000,1.5401,1.5401,1.54,1.54
20101227,191100,1.54,1.54,1.5399,1.5399
20101227,191200,1.5399,1.5399,1.5398,1.5398
20101227,191300,1.5397,1.5397,1.5397,1.5397
20101227,191400,1.5397,1.5402,1.5397,1.5402
20101227,191500,1.5403,1.5405,1.5403,1.5405
20101227,191600,1.5404,1.5404,1.5403,1.5404
20101227,191700,1.5404,1.5404,1.5401,1.5401
20101227,191800,1.5401,1.5401,1.54,1.5401
20101227,191900,1.5401,1.5401,1.5399,1.5399
20101227,192000,1.5399,1.54,1.5399,1.54
20101227,192100,1.5401,1.5401,1.5399,1.5399
20101227,192200,1.5398,1.5398,1.5397,1.5398
20101227,192300,1.5397,1.5398,1.5397,1.5398
20101227,192400,1.5398,1.5398,1.5397,1.5397
20101227,192500,1.5397,1.5398,1.5397,1.5398
20101227,192600,1.5398,1.54,1.5397,1.54
20101227,192700,1.5401,1.5401,1.5399,1.54
20101227,192800,1.54,1.54,1.54,1.54
20101227,192900,1.54,1.54,1.54,1.54
20101227,193000,1.54,1.54,1.54,1.54
20101227,193100,1.54,1.5401,1.54,1.5401
20101227,193200,1.5402,1.5403,1.5402,1.5403
20101227,193300,1.5402,1.5402,1.5401,1.5401
20101227,193400,1.5401,1.5402,1.5399,1.5399
20101227,193500,1.54,1.54,1.5399,1.54
20101227,193600,1.5401,1.5402,1.5401,1.5402
20101227,193700,1.5402,1.5402,1.5401,1.5402
20101227,193800,1.5401,1.5402,1.5401,1.5402
20101227,193900,1.5402,1.5402,1.5402,1.5402
20101227,194000,1.5402,1.5402,1.5402,1.5402
20101227,194100,1.5403,1.5403,1.5403,1.5403
20101227,194200,1.5403,1.5404,1.5403,1.5404
20101227,194300,1.5404,1.5406,1.5404,1.5405
20101227,194400,1.5406,1.5406,1.5405,1.5405
20101227,194500,1.5405,1.5405,1.5404,1.5404
20101227,194600,1.5405,1.5406,1.5405,1.5405
20101227,194700,1.5405,1.5405,1.5404,1.5404
20101227,194800,1.5404,1.5405,1.5404,1.5405
20101227,194900,1.5405,1.5406,1.5404,1.5406
20101227,195000,1.5405,1.5406,1.5405,1.5405
20101227,195100,1.5406,1.5406,1.5405,1.5405
20101227,195200,1.5405,1.5405,1.5403,1.5404
20101227,195300,1.5404,1.5405,1.5404,1.5405
20101227,195400,1.5406,1.5406,1.5402,1.5402
20101227,195500,1.5403,1.5403,1.5403,1.5403
20101227,195600,1.5403,1.5403,1.5401,1.5401
20101227,195700,1.5401,1.5401,1.54,1.54
20101227,195800,1.54,1.5401,1.54,1.54
20101227,195900,1.54,1.5402,1.54,1.5402
20101227,200000,1.5402,1.5402,1.5401,1.5402
20101227,200100,1.5402,1.5402,1.5401,1.5402
20101227,200200,1.5401,1.5402,1.5401,1.5401
20101227,200300,1.54,1.54,1.54,1.54
20101227,200400,1.54,1.54,1.54,1.54
20101227,200500,1.54,1.5401,1.54,1.5401
20101227,200600,1.54,1.5402,1.54,1.5402
20101227,200700,1.5402,1.5402,1.5402,1.5402
20101227,200800,1.5402,1.5402,1.5402,1.5402
20101227,200900,1.5402,1.5402,1.5402,1.5402
20101227,201000,1.5402,1.5402,1.5401,1.5401
20101227,201100,1.5401,1.5402,1.5401,1.5402
20101227,201200,1.5402,1.5402,1.5402,1.5402
20101227,201300,1.5401,1.5403,1.5401,1.5403
20101227,201400,1.5404,1.5406,1.5404,1.5404
20101227,201500,1.5405,1.5407,1.5405,1.5405
20101227,201600,1.5405,1.5405,1.5403,1.5403
20101227,201700,1.5402,1.5402,1.5402,1.5402
20101227,201800,1.5402,1.5402,1.5402,1.5402
20101227,201900,1.5402,1.5402,1.5402,1.5402
20101227,202000,1.5402,1.5402,1.5402,1.5402
20101227,202100,1.5402,1.5402,1.5402,1.5402
20101227,202200,1.5402,1.5404,1.5402,1.5404
20101227,202300,1.5404,1.5404,1.5404,1.5404
20101227,202400,1.5404,1.5404,1.5404,1.5404
20101227,202500,1.5404,1.5406,1.5404,1.5406
20101227,202600,1.5406,1.5407,1.5405,1.5406
20101227,202700,1.5407,1.5407,1.5406,1.5407
20101227,202800,1.5406,1.5406,1.5405,1.5405
20101227,202900,1.5406,1.5407,1.5406,1.5407
20101227,203000,1.5407,1.5407,1.5406,1.5407
20101227,203100,1.5406,1.5409,1.5406,1.5408
20101227,203200,1.5407,1.5407,1.5406,1.5406
20101227,203300,1.5406,1.5407,1.5406,1.5407
20101227,203400,1.5406,1.5406,1.5405,1.5405
20101227,203500,1.5406,1.5406,1.5405,1.5405
20101227,203600,1.5405,1.5405,1.5404,1.5405
20101227,203700,1.5405,1.5405,1.5405,1.5405
20101227,203800,1.5405,1.5406,1.5405,1.5406
20101227,203900,1.5405,1.5407,1.5405,1.5406
20101227,204000,1.5405,1.5405,1.5405,1.5405
20101227,204100,1.5405,1.5405,1.5403,1.5403
20101227,204200,1.5403,1.5404,1.5403,1.5403
20101227,204300,1.5403,1.5404,1.5403,1.5403
20101227,204400,1.5404,1.5404,1.5403,1.5403
20101227,204500,1.5404,1.5406,1.5403,1.5406
20101227,204600,1.5405,1.5405,1.5404,1.5404
20101227,204700,1.5405,1.5405,1.5403,1.5403
20101227,204800,1.5404,1.5407,1.5404,1.5407
20101227,204900,1.5406,1.5406,1.5406,1.5406
20101227,205000,1.5406,1.5406,1.5406,1.5406
20101227,205100,1.5406,1.5407,1.5406,1.5407
20101227,205200,1.5407,1.5407,1.5406,1.5406
20101227,205300,1.5407,1.5407,1.5406,1.5406
20101227,205400,1.5407,1.541,1.5406,1.5409
20101227,205500,1.5409,1.5409,1.5409,1.5409
20101227,205600,1.5408,1.5409,1.5407,1.5407
20101227,205700,1.5408,1.5408,1.5407,1.5408
20101227,205800,1.5408,1.5408,1.5408,1.5408
20101227,205900,1.5408,1.5409,1.5408,1.5408
20101227,210000,1.5409,1.5409,1.5409,1.5409
20101227,210100,1.5408,1.5413,1.5408,1.541
20101227,210200,1.5411,1.5414,1.5411,1.5414
20101227,210300,1.5413,1.5414,1.5413,1.5413
20101227,210400,1.5414,1.5416,1.5407,1.5411
20101227,210500,1.5412,1.5417,1.5411,1.5415
20101227,210600,1.5415,1.5416,1.5414,1.5415
20101227,210700,1.5415,1.5416,1.5415,1.5415
20101227,210800,1.5415,1.5416,1.5415,1.5416
20101227,210900,1.5416,1.5417,1.5416,1.5417
20101227,211000,1.5418,1.5418,1.5417,1.5418
20101227,211100,1.5417,1.5417,1.5416,1.5417
20101227,211200,1.5417,1.5417,1.5415,1.5415
20101227,211300,1.5415,1.5416,1.5415,1.5416
20101227,211400,1.5416,1.5417,1.5415,1.5417
20101227,211500,1.5418,1.5418,1.5418,1.5418
20101227,211600,1.5418,1.5418,1.5416,1.5417
20101227,211700,1.5417,1.5417,1.5417,1.5417
20101227,211800,1.5417,1.5417,1.5417,1.5417
20101227,211900,1.5417,1.5417,1.5417,1.5417
20101227,212000,1.5418,1.5418,1.5417,1.5417
20101227,212100,1.5416,1.5416,1.5415,1.5416
20101227,212200,1.5416,1.5416,1.5415,1.5416
20101227,212300,1.5416,1.5417,1.5416,1.5417
20101227,212400,1.5417,1.5417,1.5415,1.5416
20101227,212500,1.5416,1.5417,1.5416,1.5416
20101227,212600,1.5417,1.5417,1.5417,1.5417
20101227,212700,1.5418,1.5418,1.5416,1.5416
20101227,212800,1.5416,1.5416,1.5416,1.5416
20101227,212900,1.5416,1.5416,1.5416,1.5416
20101227,213000,1.5416,1.5416,1.5415,1.5416
20101227,213100,1.5416,1.5417,1.5416,1.5417
20101227,213200,1.5418,1.5418,1.5417,1.5418
20101227,213300,1.5418,1.5418,1.5418,1.5418
20101227,213400,1.5418,1.5418,1.5418,1.5418
20101227,213500,1.5418,1.5419,1.5417,1.5417
20101227,213600,1.5417,1.5417,1.5417,1.5417
20101227,213700,1.5417,1.5417,1.5417,1.5417
20101227,213800,1.5418,1.5419,1.5418,1.5418
20101227,213900,1.5417,1.5417,1.5416,1.5416
20101227,214000,1.5417,1.5418,1.5416,1.5417
20101227,214100,1.5416,1.5416,1.5416,1.5416
20101227,214200,1.5416,1.5417,1.5416,1.5416
20101227,214300,1.5416,1.5416,1.5416,1.5416
20101227,214400,1.5416,1.5417,1.5416,1.5417
20101227,214500,1.5417,1.5417,1.5417,1.5417
20101227,214600,1.5418,1.5418,1.5418,1.5418
20101227,214700,1.5418,1.5418,1.5417,1.5418
20101227,214800,1.5418,1.5418,1.5418,1.5418
20101227,214900,1.5418,1.5418,1.5418,1.5418
20101227,215000,1.5417,1.5418,1.5417,1.5418
20101227,215100,1.5418,1.5418,1.5418,1.5418
20101227,215200,1.5419,1.5419,1.5417,1.5419
20101227,215300,1.5419,1.5419,1.5419,1.5419
20101227,215400,1.5419,1.5419,1.5418,1.5418
20101227,215500,1.5418,1.5419,1.5418,1.5419
20101227,215600,1.5419,1.5419,1.5418,1.5419
20101227,215700,1.5419,1.5419,1.5418,1.5418
20101227,215800,1.5419,1.5419,1.5418,1.5418
20101227,215900,1.5419,1.5419,1.5419,1.5419
20101227,220000,1.5419,1.5419,1.5418,1.5419
20101227,220100,1.5419,1.5419,1.5419,1.5419
20101227,220200,1.5419,1.5419,1.5419,1.5419
20101227,220300,1.5419,1.5419,1.5419,1.5419
20101227,220400,1.5419,1.542,1.5419,1.542
20101227,220500,1.542,1.542,1.542,1.542
20101227,220600,1.542,1.542,1.5419,1.5419
20101227,220700,1.5419,1.542,1.5419,1.542
20101227,220800,1.542,1.542,1.542,1.542
20101227,220900,1.542,1.542,1.5419,1.5419
20101227,221000,1.5419,1.5419,1.5418,1.5419
20101227,221100,1.5419,1.542,1.5419,1.5419
20101227,221200,1.5419,1.5419,1.5419,1.5419
20101227,221300,1.5419,1.5419,1.5419,1.5419
20101227,221400,1.5419,1.5421,1.5419,1.5421
20101227,221500,1.5421,1.5421,1.5421,1.5421
20101227,221600,1.5422,1.5422,1.5421,1.5421
20101227,221700,1.5421,1.5422,1.5421,1.5421
20101227,221800,1.5421,1.5422,1.542,1.542
20101227,221900,1.542,1.542,1.542,1.542
20101227,222000,1.5419,1.5422,1.5419,1.5422
20101227,222100,1.5422,1.5422,1.5422,1.5422
20101227,222200,1.5422,1.5423,1.5422,1.5423
20101227,222300,1.5423,1.5423,1.5423,1.5423
20101227,222400,1.5422,1.5423,1.5422,1.5423
20101227,222500,1.5423,1.5423,1.5422,1.5422
20101227,222600,1.5423,1.5423,1.5423,1.5423
20101227,222700,1.5423,1.5423,1.542,1.542
20101227,222800,1.5419,1.5422,1.5419,1.5422
20101227,222900,1.5422,1.5422,1.5422,1.5422
20101227,223000,1.5422,1.5422,1.5422,1.5422
20101227,223100,1.5422,1.5422,1.5422,1.5422
20101227,223200,1.5422,1.5423,1.5422,1.5423
20101227,223300,1.5424,1.5424,1.5423,1.5423
20101227,223400,1.5424,1.5424,1.5423,1.5423
20101227,223500,1.5424,1.5425,1.5423,1.5425
20101227,223600,1.5425,1.5425,1.5425,1.5425
20101227,223700,1.5425,1.5425,1.5424,1.5424
20101227,223800,1.5424,1.5424,1.5423,1.5423
20101227,223900,1.5422,1.5423,1.5421,1.5423
20101227,224000,1.5424,1.5424,1.5424,1.5424
20101227,224100,1.5423,1.5424,1.5423,1.5424
20101227,224200,1.5424,1.5424,1.5422,1.5422
20101227,224300,1.5422,1.5422,1.5421,1.5421
20101227,224400,1.5421,1.5421,1.5421,1.5421
20101227,224500,1.542,1.542,1.542,1.542
20101227,224600,1.542,1.5421,1.542,1.5421
20101227,224700,1.5421,1.5421,1.542,1.542
20101227,224800,1.542,1.542,1.542,1.542
20101227,224900,1.542,1.542,1.542,1.542
20101227,225000,1.542,1.542,1.5419,1.5419
20101227,225100,1.5419,1.5419,1.5418,1.5419
20101227,225200,1.5418,1.5418,1.5418,1.5418
20101227,225300,1.5418,1.5418,1.5418,1.5418
20101227,225400,1.5418,1.5418,1.5418,1.5418
20101227,225500,1.5417,1.5417,1.5417,1.5417
20101227,225700,1.5416,1.5416,1.5416,1.5416
20101227,225800,1.5416,1.5416,1.5416,1.5416
20101227,230000,1.5414,1.5414,1.5414,1.5414
20101227,230200,1.5414,1.5415,1.5414,1.5415
20101227,230300,1.5414,1.5414,1.5414,1.5414
20101227,230400,1.5414,1.5415,1.5414,1.5414
20101227,230500,1.5415,1.5415,1.5415,1.5415
20101227,230600,1.5414,1.5414,1.5414,1.5414
20101227,230800,1.5414,1.5414,1.5414,1.5414
20101227,230900,1.5414,1.5415,1.5414,1.5415
20101227,231000,1.5415,1.5416,1.5415,1.5416
20101227,231100,1.5416,1.5416,1.5416,1.5416
20101227,231200,1.5416,1.5416,1.5416,1.5416
20101227,231300,1.5416,1.5417,1.5416,1.5416
20101227,231400,1.5416,1.5417,1.5416,1.5417
20101227,231500,1.5417,1.5417,1.5417,1.5417
20101227,231600,1.5419,1.5419,1.5419,1.5419
20101227,231800,1.5419,1.5419,1.5419,1.5419
20101227,231900,1.5419,1.5419,1.5419,1.5419
20101227,232000,1.5419,1.542,1.5419,1.542
20101227,232100,1.542,1.542,1.542,1.542
20101227,232200,1.542,1.542,1.542,1.542
20101227,232400,1.542,1.542,1.542,1.542
20101227,232600,1.5422,1.5422,1.5422,1.5422
20101227,232800,1.5422,1.5422,1.5422,1.5422
20101227,232900,1.5422,1.5422,1.5422,1.5422
20101227,233000,1.5425,1.5425,1.5425,1.5425
20101227,233200,1.5425,1.5425,1.5424,1.5424
20101227,233300,1.5425,1.5425,1.5425,1.5425
20101227,233400,1.5424,1.5424,1.5424,1.5424
20101227,233500,1.5424,1.5424,1.5424,1.5424
20101227,233700,1.5424,1.5424,1.5424,1.5424
20101227,233800,1.5425,1.5425,1.5424,1.5424
20101227,233900,1.5424,1.5427,1.5424,1.5427
20101227,234000,1.5427,1.5427,1.5427,1.5427
20101227,234100,1.5427,1.5427,1.5427,1.5427
20101227,234200,1.5427,1.5427,1.5427,1.5427
20101227,234400,1.5427,1.5427,1.5427,1.5427
20101227,234500,1.5427,1.5427,1.5427,1.5427
20101227,234600,1.5427,1.5427,1.5427,1.5427
20101227,234700,1.5433,1.5433,1.5433,1.5433
20101227,234900,1.5433,1.5433,1.5433,1.5433
20101227,235000,1.5434,1.5434,1.5434,1.5434
20101227,235200,1.5434,1.5434,1.5434,1.5434
20101227,235300,1.5433,1.5434,1.5433,1.5433
20101227,235400,1.5436,1.5436,1.5436,1.5436
20101227,235600,1.5439,1.5439,1.5439,1.5439
20101227,235800,1.5439,1.544,1.5439,1.544
20101227,235900,1.5439,1.544,1.5438,1.5439
20101228,0,1.544,1.544,1.544,1.544
20101228,100,1.5442,1.5442,1.5442,1.5442
20101228,200,1.5441,1.5441,1.5441,1.5441
20101228,400,1.5441,1.5441,1.5441,1.5441
20101228,500,1.5442,1.5442,1.5442,1.5442
20101228,600,1.5442,1.5442,1.5442,1.5442
20101228,700,1.5446,1.5446,1.5446,1.5446
20101228,900,1.5445,1.5445,1.5444,1.5444
20101228,1000,1.5445,1.5445,1.5445,1.5445
20101228,1100,1.5443,1.5443,1.5443,1.5443
20101228,1200,1.5445,1.5445,1.5445,1.5445
20101228,1400,1.5452,1.5452,1.5452,1.5452
20101228,1600,1.547,1.547,1.547,1.547
20101228,1700,1.5472,1.5472,1.5472,1.5472
20101228,1800,1.5463,1.5463,1.5463,1.5463
20101228,1900,1.5467,1.5467,1.5467,1.5467
20101228,2000,1.5474,1.5474,1.5474,1.5474
20101228,2100,1.5472,1.5472,1.5472,1.5472
20101228,2200,1.5472,1.5472,1.5472,1.5472
20101228,2300,1.5472,1.5472,1.5472,1.5472
20101228,2400,1.5471,1.5471,1.5471,1.5471
20101228,2500,1.5475,1.5475,1.5475,1.5475
20101228,2600,1.5474,1.5474,1.5474,1.5474
20101228,2700,1.5476,1.5476,1.5476,1.5476
20101228,2900,1.5476,1.5476,1.5476,1.5476
20101228,3000,1.5484,1.5484,1.5484,1.5484
20101228,3100,1.5472,1.5472,1.5472,1.5472
20101228,3200,1.5474,1.5474,1.5474,1.5474
20101228,3400,1.5473,1.5475,1.5471,1.5473
20101228,3500,1.5472,1.5472,1.5472,1.5472
20101228,3600,1.5473,1.5473,1.5473,1.5473
20101228,3700,1.5471,1.5471,1.5471,1.5471
20101228,3800,1.5471,1.5471,1.5471,1.5471
20101228,3900,1.5472,1.5472,1.5472,1.5472
20101228,4000,1.5471,1.5471,1.5471,1.5471
20101228,4200,1.5471,1.5472,1.5471,1.5471
20101228,4300,1.5471,1.5474,1.5471,1.5474
20101228,4400,1.5475,1.5475,1.5473,1.5473
20101228,4500,1.5477,1.5477,1.5477,1.5477
20101228,4700,1.5476,1.5477,1.5476,1.5476
20101228,4800,1.5476,1.5476,1.5475,1.5475
20101228,4900,1.5476,1.5476,1.5475,1.5476
20101228,5000,1.5479,1.5479,1.5479,1.5479
20101228,5100,1.5481,1.5481,1.5481,1.5481
20101228,5200,1.5481,1.5481,1.5481,1.5481
20101228,5400,1.5472,1.5472,1.5472,1.5472
20101228,5500,1.5473,1.5473,1.5473,1.5473
20101228,5700,1.547,1.547,1.547,1.547
20101228,5900,1.5471,1.5471,1.547,1.5471
20101228,10000,1.547,1.547,1.547,1.547
20101228,10100,1.547,1.547,1.547,1.547
20101228,10400,1.547,1.547,1.547,1.547
20101228,10500,1.5469,1.5469,1.5469,1.5469
20101228,10600,1.5471,1.5471,1.5471,1.5471
20101228,10800,1.547,1.547,1.547,1.547
20101228,10900,1.5467,1.5467,1.5467,1.5467
20101228,11000,1.5469,1.5469,1.5469,1.5469
20101228,11100,1.5469,1.5469,1.5469,1.5469
20101228,11200,1.5469,1.5469,1.5469,1.5469
20101228,11400,1.5476,1.5476,1.5476,1.5476
20101228,11500,1.5474,1.5474,1.5474,1.5474
20101228,11600,1.5471,1.5471,1.5471,1.5471
20101228,11700,1.5471,1.5471,1.5471,1.5471
20101228,11800,1.5473,1.5473,1.5473,1.5473
20101228,12000,1.5473,1.5475,1.5472,1.5475
20101228,12100,1.5475,1.5475,1.5472,1.5473
20101228,12200,1.5473,1.5473,1.5472,1.5472
20101228,12300,1.5471,1.5472,1.5471,1.5472
20101228,12400,1.5472,1.5474,1.5472,1.5474
20101228,12500,1.5474,1.5474,1.5474,1.5474
20101228,12700,1.5474,1.5474,1.5474,1.5474
20101228,12800,1.5472,1.5472,1.5472,1.5472
20101228,12900,1.5472,1.5472,1.5472,1.5472
20101228,13000,1.5473,1.5473,1.5473,1.5473
20101228,13100,1.5474,1.5474,1.5474,1.5474
20101228,13200,1.5474,1.5474,1.5474,1.5474
20101228,13300,1.5474,1.5474,1.5474,1.5474
20101228,13500,1.5469,1.5469,1.5469,1.5469
20101228,13600,1.5469,1.5469,1.5469,1.5469
20101228,13700,1.5469,1.5469,1.5469,1.5469
20101228,13800,1.5468,1.5468,1.5468,1.5468
20101228,13900,1.5468,1.5468,1.5468,1.5468
20101228,14100,1.5468,1.5468,1.5466,1.5466
20101228,14200,1.5466,1.5466,1.5466,1.5466
20101228,14300,1.5466,1.5466,1.5466,1.5466
20101228,14500,1.5469,1.5469,1.5469,1.5469
20101228,14700,1.5469,1.5469,1.5469,1.5469
20101228,14900,1.5469,1.5469,1.5467,1.5469
20101228,15000,1.5468,1.5469,1.5468,1.5468
20101228,15100,1.5469,1.5469,1.5467,1.5467
20101228,15200,1.5467,1.5467,1.5467,1.5467
20101228,15300,1.5469,1.5469,1.5469,1.5469
20101228,15400,1.5466,1.5466,1.5466,1.5466
20101228,15500,1.5467,1.5467,1.5467,1.5467
20101228,15700,1.5466,1.5466,1.5466,1.5466
20101228,15800,1.5466,1.5467,1.5466,1.5466
20101228,15900,1.5466,1.5466,1.5466,1.5466
20101228,20000,1.5466,1.5466,1.5466,1.5466
20101228,20200,1.5467,1.5467,1.5467,1.5467
20101228,20400,1.5466,1.5466,1.5466,1.5466
20101228,20500,1.5466,1.5466,1.5466,1.5466
20101228,20600,1.5467,1.5467,1.5467,1.5467
20101228,20800,1.5466,1.5466,1.5466,1.5466
20101228,21000,1.5468,1.5468,1.5468,1.5468
20101228,21200,1.5467,1.5468,1.5467,1.5467
20101228,21300,1.5466,1.5466,1.5466,1.5466
20101228,21500,1.5467,1.5467,1.5467,1.5467
20101228,21600,1.5468,1.5468,1.5468,1.5468
20101228,21800,1.5468,1.5468,1.5468,1.5468
20101228,21900,1.5468,1.5468,1.5468,1.5468
20101228,22000,1.5468,1.5468,1.5468,1.5468
20101228,22100,1.5468,1.5468,1.5468,1.5468
20101228,22200,1.5468,1.5468,1.5468,1.5468
20101228,22300,1.5467,1.5467,1.5467,1.5467
20101228,22400,1.5466,1.5466,1.5466,1.5466
20101228,22600,1.5466,1.5468,1.5466,1.5468
20101228,22700,1.5468,1.5468,1.5468,1.5468
20101228,22800,1.5468,1.5468,1.5468,1.5468
20101228,22900,1.5466,1.5466,1.5466,1.5466
20101228,23000,1.5466,1.5466,1.5466,1.5466
20101228,23200,1.5467,1.5467,1.5466,1.5467
20101228,23300,1.547,1.547,1.547,1.547
20101228,23500,1.547,1.547,1.547,1.547
20101228,23600,1.547,1.5471,1.547,1.5471
20101228,23700,1.5473,1.5473,1.5473,1.5473
20101228,23900,1.5472,1.5472,1.5472,1.5472
20101228,24100,1.5474,1.5474,1.5474,1.5474
20101228,24200,1.5473,1.5473,1.5473,1.5473
20101228,24300,1.547,1.547,1.547,1.547
20101228,24400,1.5471,1.5471,1.5471,1.5471
20101228,24500,1.5469,1.5469,1.5469,1.5469
20101228,24600,1.5469,1.5469,1.5469,1.5469
20101228,24800,1.5469,1.5469,1.5469,1.5469
20101228,24900,1.547,1.547,1.547,1.547
20101228,25000,1.5469,1.5469,1.5469,1.5469
20101228,25100,1.5468,1.5468,1.5468,1.5468
20101228,25300,1.5469,1.5469,1.5469,1.5469
20101228,25400,1.547,1.547,1.547,1.547
20101228,25600,1.5466,1.5466,1.5466,1.5466
20101228,25700,1.5466,1.5466,1.5466,1.5466
20101228,25900,1.5467,1.5467,1.5467,1.5467
20101228,30100,1.5468,1.5468,1.5468,1.5468
20101228,30300,1.5469,1.5469,1.5469,1.5469
20101228,30400,1.5469,1.5469,1.5469,1.5469
20101228,30500,1.547,1.547,1.547,1.547
20101228,30700,1.547,1.547,1.5467,1.5468
20101228,30800,1.5469,1.5469,1.5469,1.5469
20101228,31000,1.5469,1.547,1.5469,1.5469
20101228,31100,1.547,1.547,1.5468,1.547
20101228,31200,1.5469,1.547,1.5469,1.547
20101228,31300,1.5471,1.5471,1.5471,1.5471
20101228,31400,1.5471,1.5471,1.547,1.5471
20101228,31500,1.5471,1.5471,1.547,1.5471
20101228,31600,1.5471,1.5471,1.547,1.547
20101228,31700,1.5471,1.5471,1.5471,1.5471
20101228,31800,1.5472,1.5473,1.547,1.547
20101228,31900,1.547,1.5471,1.547,1.547
20101228,32000,1.547,1.547,1.5469,1.5469
20101228,32100,1.5469,1.5469,1.5469,1.5469
20101228,32200,1.5469,1.5469,1.5469,1.5469
20101228,32300,1.5469,1.5469,1.5469,1.5469
20101228,32500,1.547,1.547,1.547,1.547
20101228,32600,1.547,1.547,1.547,1.547
20101228,32700,1.547,1.547,1.547,1.547
20101228,32800,1.547,1.547,1.547,1.547
20101228,33000,1.5469,1.547,1.5468,1.5469
20101228,33100,1.5469,1.5469,1.5469,1.5469
20101228,33200,1.5469,1.5469,1.5469,1.5469
20101228,33300,1.5469,1.5469,1.5467,1.5467
20101228,33400,1.5468,1.5469,1.5468,1.5469
20101228,33500,1.547,1.5472,1.547,1.5471
20101228,33600,1.5472,1.5472,1.5472,1.5472
20101228,33700,1.5472,1.5472,1.5472,1.5472
20101228,33800,1.5474,1.5474,1.5474,1.5474
20101228,34000,1.5474,1.5474,1.5473,1.5473
20101228,34100,1.5474,1.5474,1.5474,1.5474
20101228,34200,1.5473,1.5473,1.5473,1.5473
20101228,34300,1.5475,1.5475,1.5475,1.5475
20101228,34400,1.5476,1.5476,1.5476,1.5476
20101228,34500,1.5476,1.5476,1.5476,1.5476
20101228,34600,1.5476,1.5476,1.5476,1.5476
20101228,34700,1.5476,1.5476,1.5476,1.5476
20101228,34800,1.5476,1.5476,1.5476,1.5476
20101228,34900,1.5475,1.5475,1.5475,1.5475
20101228,35100,1.5475,1.5475,1.5473,1.5473
20101228,35200,1.5472,1.5473,1.5472,1.5472
20101228,35300,1.5472,1.5472,1.5471,1.5472
20101228,35400,1.5472,1.5472,1.5471,1.5472
20101228,35500,1.5471,1.5473,1.5471,1.5473
20101228,35600,1.5472,1.5475,1.5471,1.5474
20101228,35700,1.548,1.548,1.548,1.548
20101228,35800,1.5481,1.5481,1.5481,1.5481
20101228,35900,1.5483,1.5483,1.5483,1.5483
20101228,40000,1.548,1.548,1.548,1.548
20101228,40200,1.548,1.548,1.5476,1.5476
20101228,40300,1.5476,1.5476,1.5476,1.5476
20101228,40400,1.5477,1.5477,1.5477,1.5477
20101228,40500,1.5477,1.5477,1.5477,1.5477
20101228,40600,1.5476,1.5476,1.5476,1.5476
20101228,40700,1.5477,1.5477,1.5477,1.5477
20101228,40800,1.5475,1.5475,1.5475,1.5475
20101228,41000,1.5476,1.5476,1.5476,1.5476
20101228,41200,1.5481,1.5481,1.5481,1.5481
20101228,41400,1.548,1.548,1.548,1.548
20101228,41600,1.5482,1.5482,1.5482,1.5482
20101228,41800,1.5482,1.5483,1.5482,1.5482
20101228,41900,1.548,1.548,1.548,1.548
20101228,42000,1.5475,1.5475,1.5475,1.5475
20101228,42200,1.5475,1.5476,1.5475,1.5475
20101228,42300,1.5471,1.5471,1.5471,1.5471
20101228,42400,1.5471,1.5471,1.5471,1.5471
20101228,42500,1.5471,1.5471,1.5471,1.5471
20101228,42600,1.5473,1.5473,1.5473,1.5473
20101228,42800,1.5473,1.5473,1.5473,1.5473
20101228,42900,1.5472,1.5473,1.5471,1.5471
20101228,43000,1.5472,1.5472,1.5472,1.5472
20101228,43100,1.5472,1.5472,1.5472,1.5472
20101228,43300,1.5472,1.5473,1.5472,1.5473
20101228,43400,1.5477,1.5477,1.5477,1.5477
20101228,43600,1.5477,1.5477,1.5477,1.5477
20101228,43800,1.5477,1.5478,1.5477,1.5477
20101228,43900,1.5477,1.5477,1.5477,1.5477
20101228,44000,1.5477,1.5479,1.5477,1.5479
20101228,44100,1.548,1.548,1.5479,1.5479
20101228,44200,1.5479,1.5479,1.5477,1.5477
20101228,44300,1.5477,1.5477,1.5477,1.5477
20101228,44400,1.5481,1.5481,1.5481,1.5481
20101228,44600,1.5482,1.5482,1.548,1.5481
20101228,44700,1.5481,1.5481,1.5481,1.5481
20101228,44800,1.5481,1.5481,1.5481,1.5481
20101228,44900,1.5481,1.5481,1.5481,1.5481
20101228,45100,1.5481,1.5482,1.5481,1.5482
20101228,45200,1.5482,1.5482,1.5482,1.5482
20101228,45400,1.5481,1.5482,1.5478,1.5479
20101228,45500,1.5479,1.5479,1.5479,1.5479
20101228,45600,1.5479,1.5479,1.5479,1.5479
20101228,45700,1.5479,1.5481,1.5479,1.5481
20101228,45800,1.5481,1.5481,1.5479,1.5479
20101228,45900,1.5479,1.548,1.5479,1.548
20101228,50000,1.548,1.5481,1.548,1.548
20101228,50100,1.5479,1.5481,1.5478,1.5481
20101228,50200,1.5481,1.5481,1.5481,1.5481
20101228,50300,1.5483,1.5483,1.5483,1.5483
20101228,50400,1.5481,1.5481,1.5481,1.5481
20101228,50500,1.548,1.548,1.548,1.548
20101228,50600,1.5482,1.5482,1.5482,1.5482
20101228,50800,1.5481,1.5481,1.5481,1.5481
20101228,51000,1.5481,1.5481,1.5481,1.5481
20101228,51100,1.548,1.548,1.548,1.548
20101228,51200,1.548,1.548,1.548,1.548
20101228,51300,1.548,1.548,1.548,1.548
20101228,51500,1.5479,1.5479,1.5479,1.5479
20101228,51600,1.548,1.548,1.548,1.548
20101228,51700,1.548,1.548,1.548,1.548
20101228,51800,1.548,1.548,1.548,1.548
20101228,52000,1.5479,1.5479,1.5479,1.5479
20101228,52200,1.5479,1.5479,1.5479,1.5479
20101228,52300,1.548,1.548,1.548,1.548
20101228,52400,1.5479,1.5479,1.5479,1.5479
20101228,52600,1.5478,1.5478,1.5478,1.5478
20101228,52700,1.5479,1.5479,1.5479,1.5479
20101228,52800,1.5481,1.5481,1.5481,1.5481
20101228,53000,1.548,1.5484,1.548,1.5484
20101228,53100,1.5483,1.5483,1.5483,1.5483
20101228,53200,1.5485,1.5485,1.5485,1.5485
20101228,53400,1.5484,1.5484,1.5484,1.5484
20101228,53500,1.5485,1.5485,1.5485,1.5485
20101228,53700,1.5485,1.5485,1.5485,1.5485
20101228,53800,1.5485,1.5485,1.5485,1.5485
20101228,53900,1.5484,1.5484,1.5484,1.5484
20101228,54000,1.5484,1.5484,1.5484,1.5484
20101228,54100,1.5483,1.5483,1.5483,1.5483
20101228,54200,1.5483,1.5483,1.5483,1.5483
20101228,54400,1.5483,1.5484,1.5483,1.5483
20101228,54500,1.5483,1.5483,1.5483,1.5483
20101228,54700,1.5483,1.5483,1.5479,1.5479
20101228,54800,1.5478,1.5478,1.5478,1.5478
20101228,55000,1.5478,1.5478,1.5477,1.5477
20101228,55100,1.5477,1.5477,1.5477,1.5477
20101228,55200,1.5475,1.5475,1.5475,1.5475
20101228,55300,1.5473,1.5473,1.5473,1.5473
20101228,55500,1.5473,1.5473,1.5473,1.5473
20101228,55600,1.5474,1.5474,1.5474,1.5474
20101228,55800,1.5474,1.5474,1.5474,1.5474
20101228,55900,1.5474,1.5474,1.5473,1.5473
20101228,60000,1.5473,1.5474,1.5473,1.5474
20101228,60100,1.5474,1.5475,1.5474,1.5474
20101228,60200,1.5475,1.5475,1.5475,1.5475
20101228,60400,1.5474,1.5474,1.5474,1.5474
20101228,60500,1.5474,1.5474,1.5474,1.5474
20101228,60600,1.5474,1.5474,1.5474,1.5474
20101228,60700,1.5474,1.5474,1.5474,1.5474
20101228,60800,1.5474,1.5474,1.5474,1.5474
20101228,61000,1.5474,1.5475,1.5473,1.5474
20101228,61100,1.5474,1.5475,1.5474,1.5474
20101228,61200,1.5475,1.5475,1.5474,1.5474
20101228,61300,1.5475,1.5476,1.5475,1.5476
20101228,61400,1.5475,1.5475,1.5475,1.5475
20101228,61500,1.5475,1.5475,1.5475,1.5475
20101228,61600,1.5474,1.5474,1.5474,1.5474
20101228,61700,1.5475,1.5475,1.5475,1.5475
20101228,61800,1.5475,1.5475,1.5475,1.5475
20101228,61900,1.5474,1.5474,1.5474,1.5474
20101228,62000,1.5466,1.5466,1.5466,1.5466
20101228,62100,1.5464,1.5464,1.5464,1.5464
20101228,62200,1.5465,1.5465,1.5465,1.5465
20101228,62300,1.5465,1.5465,1.5465,1.5465
20101228,62400,1.5465,1.5465,1.5465,1.5465
20101228,62600,1.5469,1.5469,1.5469,1.5469
20101228,62800,1.5469,1.5469,1.5469,1.5469
20101228,62900,1.5469,1.5469,1.5469,1.5469
20101228,63000,1.5469,1.5469,1.5469,1.5469
20101228,63200,1.5469,1.5469,1.5467,1.5467
20101228,63300,1.5468,1.5468,1.5467,1.5467
20101228,63400,1.5467,1.5467,1.5465,1.5465
20101228,63500,1.5465,1.5466,1.5465,1.5465
20101228,63600,1.5464,1.5464,1.5464,1.5464
20101228,63700,1.5463,1.5463,1.5463,1.5463
20101228,63800,1.5464,1.5464,1.5464,1.5464
20101228,64000,1.5464,1.5464,1.5464,1.5464
20101228,64100,1.5464,1.5464,1.5464,1.5464
20101228,64200,1.5463,1.5463,1.5463,1.5463
20101228,64300,1.5463,1.5463,1.5463,1.5463
20101228,64500,1.5463,1.5463,1.5462,1.5462
20101228,64600,1.5462,1.5462,1.5461,1.5462
20101228,64700,1.5462,1.5462,1.5462,1.5462
20101228,64800,1.5462,1.5462,1.5461,1.5461
20101228,64900,1.5462,1.5467,1.5461,1.5467
20101228,65000,1.5466,1.5466,1.5464,1.5465
20101228,65100,1.5463,1.5463,1.5463,1.5463
20101228,65300,1.5463,1.5464,1.5463,1.5463
20101228,65400,1.5464,1.5464,1.5463,1.5463
20101228,65500,1.5464,1.5466,1.5464,1.5466
20101228,65600,1.5466,1.5467,1.5466,1.5466
20101228,65700,1.5462,1.5462,1.5462,1.5462
20101228,65800,1.5462,1.5462,1.5462,1.5462
20101228,70000,1.5458,1.5458,1.5458,1.5458
20101228,70100,1.546,1.546,1.546,1.546
20101228,70200,1.5463,1.5463,1.5463,1.5463
20101228,70300,1.5464,1.5464,1.5464,1.5464
20101228,70500,1.5468,1.5468,1.5468,1.5468
20101228,70700,1.5469,1.5469,1.5468,1.5468
20101228,70800,1.5469,1.5469,1.5469,1.5469
20101228,70900,1.5469,1.5469,1.5469,1.5469
20101228,71100,1.5468,1.5468,1.5468,1.5468
20101228,71300,1.5468,1.5468,1.5467,1.5468
20101228,71400,1.5468,1.5469,1.5468,1.5469
20101228,71500,1.5471,1.5471,1.5471,1.5471
20101228,71600,1.5471,1.5471,1.5471,1.5471
20101228,71800,1.5471,1.5471,1.5471,1.5471
20101228,71900,1.5472,1.5472,1.5472,1.5472
20101228,72000,1.5467,1.5467,1.5467,1.5467
20101228,72100,1.5467,1.5467,1.5467,1.5467
20101228,72200,1.5465,1.5465,1.5465,1.5465
20101228,72400,1.5466,1.5466,1.5465,1.5466
20101228,72500,1.5465,1.5465,1.5462,1.5462
20101228,72600,1.5462,1.5463,1.5462,1.5463
20101228,72700,1.5464,1.5467,1.5464,1.5466
20101228,72800,1.5466,1.5466,1.5466,1.5466
20101228,72900,1.5466,1.5466,1.5466,1.5466
20101228,73100,1.5467,1.5467,1.5464,1.5464
20101228,73200,1.5463,1.5464,1.5462,1.5463
20101228,73300,1.5462,1.5464,1.5462,1.5464
20101228,73400,1.5464,1.5464,1.5463,1.5464
20101228,73500,1.5464,1.5464,1.5464,1.5464
20101228,73700,1.5463,1.5464,1.5462,1.5464
20101228,73800,1.5464,1.5464,1.5464,1.5464
20101228,74000,1.546,1.546,1.546,1.546
20101228,74100,1.5458,1.5458,1.5458,1.5458
20101228,74200,1.5458,1.5458,1.5458,1.5458
20101228,74400,1.5458,1.5458,1.5458,1.5458
20101228,74500,1.5458,1.5458,1.5458,1.5458
20101228,74700,1.5457,1.5458,1.5457,1.5457
20101228,74800,1.5458,1.5458,1.5457,1.5457
20101228,74900,1.543,1.543,1.543,1.543
20101228,75100,1.5435,1.5435,1.5435,1.5435
20101228,75300,1.5434,1.5435,1.5434,1.5434
20101228,75400,1.5435,1.5435,1.5435,1.5435
20101228,75500,1.5435,1.5435,1.5435,1.5435
20101228,75700,1.5436,1.5436,1.5436,1.5436
20101228,75800,1.5432,1.5432,1.5432,1.5432
20101228,75900,1.5429,1.5429,1.5429,1.5429
20101228,80000,1.5429,1.5429,1.5429,1.5429
20101228,80100,1.5426,1.5426,1.5426,1.5426
20101228,80300,1.5429,1.5429,1.5429,1.5429
20101228,80500,1.5435,1.5435,1.5435,1.5435
20101228,80600,1.5434,1.5434,1.5434,1.5434
20101228,80700,1.5439,1.5439,1.5439,1.5439
20101228,80900,1.5439,1.5439,1.5439,1.5439
20101228,81000,1.5441,1.5441,1.5441,1.5441
20101228,81100,1.5442,1.5442,1.5442,1.5442
20101228,81200,1.5442,1.5442,1.5442,1.5442
20101228,81300,1.5442,1.5442,1.5442,1.5442
20101228,81500,1.5442,1.5443,1.5442,1.5443
20101228,81600,1.5442,1.5442,1.5442,1.5442
20101228,81700,1.5442,1.5442,1.5442,1.5442
20101228,81800,1.5443,1.5443,1.5443,1.5443
20101228,81900,1.5444,1.5444,1.5444,1.5444
20101228,82000,1.5444,1.5444,1.5444,1.5444
20101228,82100,1.5445,1.5445,1.5445,1.5445
20101228,82200,1.5444,1.5444,1.5444,1.5444
20101228,82400,1.5444,1.5444,1.5444,1.5444
20101228,82600,1.544,1.544,1.544,1.544
20101228,82700,1.5442,1.5442,1.5442,1.5442
20101228,82900,1.5441,1.5441,1.5441,1.5441
20101228,83100,1.5442,1.5442,1.544,1.544
20101228,83200,1.5442,1.5442,1.5442,1.5442
20101228,83400,1.5442,1.5443,1.5441,1.5442
20101228,83500,1.5441,1.5441,1.544,1.5441
20101228,83600,1.544,1.5441,1.5439,1.5439
20101228,83700,1.5439,1.5439,1.5439,1.5439
20101228,83800,1.5443,1.5443,1.5443,1.5443
20101228,84000,1.544,1.544,1.544,1.544
20101228,84100,1.5445,1.5445,1.5445,1.5445
20101228,84300,1.5444,1.5444,1.5441,1.5442
20101228,84400,1.544,1.544,1.544,1.544
20101228,84500,1.5446,1.5446,1.5446,1.5446
20101228,84600,1.5441,1.5441,1.5441,1.5441
20101228,84700,1.5437,1.5437,1.5437,1.5437
20101228,84800,1.5436,1.5436,1.5436,1.5436
20101228,84900,1.544,1.544,1.544,1.544
20101228,85100,1.5439,1.5442,1.5439,1.5442
20101228,85200,1.5443,1.5443,1.5443,1.5443
20101228,85300,1.5444,1.5444,1.5444,1.5444
20101228,85500,1.5443,1.5445,1.5442,1.5445
20101228,85600,1.5445,1.5445,1.5445,1.5445
20101228,85700,1.5446,1.5446,1.5446,1.5446
20101228,85900,1.5445,1.5445,1.5445,1.5445
20101228,90000,1.5443,1.5443,1.5443,1.5443
20101228,90200,1.544,1.544,1.544,1.544
20101228,90400,1.544,1.544,1.5438,1.5438
20101228,90500,1.5438,1.5438,1.5438,1.5438
20101228,90600,1.5437,1.5437,1.5437,1.5437
20101228,90800,1.5437,1.5437,1.5436,1.5436
20101228,90900,1.5437,1.5438,1.5437,1.5438
20101228,91000,1.5439,1.5439,1.5439,1.5439
20101228,91100,1.5439,1.5439,1.5439,1.5439
20101228,91300,1.5438,1.5439,1.5438,1.5439
20101228,91400,1.544,1.544,1.544,1.544
20101228,91600,1.544,1.544,1.5439,1.544
20101228,91700,1.5441,1.5441,1.544,1.5441
20101228,91800,1.5441,1.5441,1.5441,1.5441
20101228,92000,1.5439,1.5439,1.5439,1.5439
20101228,92100,1.5439,1.5439,1.5439,1.5439
20101228,92300,1.5438,1.5439,1.5438,1.5439
20101228,92400,1.5438,1.5438,1.5438,1.5438
20101228,92500,1.5438,1.5439,1.5437,1.5438
20101228,92600,1.5437,1.5437,1.5437,1.5437
20101228,92800,1.5436,1.5437,1.5435,1.5435
20101228,92900,1.5434,1.5434,1.5434,1.5434
20101228,93000,1.5433,1.5433,1.5433,1.5433
20101228,93200,1.5432,1.5432,1.5432,1.5432
20101228,93300,1.5432,1.5432,1.5432,1.5432
20101228,93400,1.543,1.543,1.543,1.543
20101228,93500,1.5431,1.5431,1.5431,1.5431
20101228,93600,1.543,1.543,1.543,1.543
20101228,93700,1.5431,1.5431,1.5431,1.5431
20101228,93800,1.543,1.543,1.543,1.543
20101228,93900,1.543,1.543,1.543,1.543
20101228,94000,1.543,1.543,1.543,1.543
20101228,94100,1.5429,1.5429,1.5429,1.5429
20101228,94300,1.5429,1.5429,1.5428,1.5428
20101228,94400,1.5429,1.5429,1.5428,1.5428
20101228,94500,1.5429,1.5429,1.5429,1.5429
20101228,94600,1.5428,1.5428,1.5428,1.5428
20101228,94800,1.5428,1.5428,1.5428,1.5428
20101228,94900,1.5416,1.5416,1.5416,1.5416
20101228,95000,1.5415,1.5415,1.5415,1.5415
20101228,95100,1.5417,1.5417,1.5417,1.5417
20101228,95200,1.5416,1.5416,1.5416,1.5416
20101228,95400,1.5415,1.5415,1.5415,1.5415
20101228,95500,1.5418,1.5418,1.5418,1.5418
20101228,95700,1.5422,1.5422,1.5422,1.5422
20101228,95800,1.5425,1.5425,1.5425,1.5425
20101228,95900,1.5432,1.5432,1.5432,1.5432
20101228,100000,1.543,1.543,1.543,1.543
20101228,100100,1.5431,1.5431,1.5431,1.5431
20101228,100200,1.543,1.543,1.543,1.543
20101228,100400,1.5431,1.5431,1.5427,1.5428
20101228,100500,1.5428,1.5429,1.5427,1.5427
20101228,100600,1.543,1.543,1.543,1.543
20101228,100800,1.5425,1.5425,1.5425,1.5425
20101228,101000,1.5424,1.5424,1.5423,1.5423
20101228,101100,1.5424,1.5424,1.5423,1.5424
20101228,101200,1.5424,1.5424,1.5423,1.5424
20101228,101300,1.5424,1.5424,1.5424,1.5424
20101228,101400,1.5426,1.5426,1.5426,1.5426
20101228,101500,1.5429,1.5429,1.5429,1.5429
20101228,101600,1.5427,1.5427,1.5427,1.5427
20101228,101700,1.5425,1.5425,1.5425,1.5425
20101228,101800,1.5426,1.5426,1.5426,1.5426
20101228,101900,1.5423,1.5423,1.5423,1.5423
20101228,102000,1.5417,1.5417,1.5417,1.5417
20101228,102200,1.5416,1.5419,1.5416,1.5417
20101228,102300,1.5417,1.5417,1.5417,1.5417
20101228,102400,1.5419,1.5419,1.5419,1.5419
20101228,102500,1.5417,1.5417,1.5417,1.5417
20101228,102700,1.5418,1.5419,1.5417,1.5418
20101228,102800,1.5419,1.5421,1.5417,1.5418
20101228,102900,1.542,1.542,1.542,1.542
20101228,103000,1.5423,1.5423,1.5423,1.5423
20101228,103200,1.5424,1.5424,1.5424,1.5424
20101228,103300,1.5425,1.5425,1.5425,1.5425
20101228,103400,1.5425,1.5425,1.5425,1.5425
20101228,103600,1.5423,1.5423,1.5423,1.5423
20101228,103800,1.5422,1.5424,1.5421,1.5424
20101228,103900,1.5422,1.5422,1.5422,1.5422
20101228,104100,1.5422,1.5423,1.5421,1.5423
20101228,104200,1.5422,1.5422,1.5418,1.5418
20101228,104300,1.5418,1.5418,1.5417,1.5418
20101228,104400,1.5418,1.5423,1.5418,1.5423
20101228,104500,1.5422,1.5423,1.5421,1.5422
20101228,104600,1.5423,1.5423,1.5423,1.5423
20101228,104800,1.5424,1.5425,1.5424,1.5424
20101228,104900,1.5423,1.5423,1.5423,1.5423
20101228,105100,1.5424,1.5424,1.5423,1.5423
20101228,105200,1.5423,1.5423,1.5423,1.5423
20101228,105400,1.5424,1.5425,1.5423,1.5425
20101228,105500,1.5425,1.5428,1.5425,1.5426
20101228,105600,1.5428,1.5428,1.5428,1.5428
20101228,105800,1.5429,1.543,1.5427,1.5427
20101228,105900,1.5419,1.5419,1.5419,1.5419
20101228,110000,1.5419,1.5419,1.5419,1.5419
20101228,110100,1.5419,1.5419,1.5419,1.5419
20101228,110200,1.5415,1.5415,1.5415,1.5415
20101228,110300,1.5411,1.5411,1.5411,1.5411
20101228,110400,1.5411,1.5411,1.5411,1.5411
20101228,110500,1.5413,1.5413,1.5413,1.5413
20101228,110600,1.542,1.542,1.542,1.542
20101228,110700,1.5422,1.5422,1.5422,1.5422
20101228,110900,1.5425,1.5425,1.5425,1.5425
20101228,111000,1.5423,1.5423,1.5423,1.5423
20101228,111200,1.5423,1.5423,1.5423,1.5423
20101228,111300,1.5423,1.5423,1.5423,1.5423
20101228,111500,1.5423,1.5424,1.5423,1.5423
20101228,111600,1.542,1.542,1.542,1.542
20101228,111700,1.5423,1.5423,1.5423,1.5423
20101228,111900,1.5425,1.5425,1.5425,1.5425
20101228,112000,1.5417,1.5417,1.5417,1.5417
20101228,112100,1.5424,1.5424,1.5424,1.5424
20101228,112300,1.5424,1.5424,1.5424,1.5424
20101228,112400,1.5425,1.5425,1.5425,1.5425
20101228,112500,1.5424,1.5424,1.5424,1.5424
20101228,112600,1.5427,1.5427,1.5427,1.5427
20101228,112800,1.5427,1.5428,1.5427,1.5428
20101228,112900,1.5433,1.5433,1.5433,1.5433
20101228,113100,1.5432,1.5436,1.543,1.5436
20101228,113200,1.5439,1.5439,1.5439,1.5439
20101228,113300,1.544,1.544,1.544,1.544
20101228,113500,1.5441,1.5447,1.5441,1.5446
20101228,113600,1.5457,1.5457,1.5457,1.5457
20101228,113700,1.5454,1.5454,1.5454,1.5454
20101228,113900,1.5455,1.5456,1.5454,1.5455
20101228,114000,1.546,1.546,1.546,1.546
20101228,114100,1.5469,1.5469,1.5469,1.5469
20101228,114300,1.5468,1.5468,1.5464,1.5466
20101228,114400,1.548,1.548,1.548,1.548
20101228,114500,1.548,1.548,1.548,1.548
20101228,114600,1.548,1.548,1.548,1.548
20101228,114800,1.548,1.548,1.5478,1.5479
20101228,114900,1.548,1.5481,1.5477,1.5477
20101228,115000,1.5479,1.5479,1.5479,1.5479
20101228,115100,1.5481,1.5481,1.5481,1.5481
20101228,115200,1.549,1.549,1.549,1.549
20101228,115300,1.5507,1.5507,1.5507,1.5507
20101228,115400,1.5505,1.5505,1.5505,1.5505
20101228,115600,1.5503,1.5503,1.5503,1.5503
20101228,115700,1.5502,1.5502,1.5502,1.5502
20101228,115800,1.5497,1.5497,1.5497,1.5497
20101228,120000,1.5503,1.5503,1.5503,1.5503
20101228,120200,1.5504,1.5504,1.55,1.55
20101228,120300,1.5498,1.5498,1.5498,1.5498
20101228,120500,1.5496,1.5496,1.5496,1.5496
20101228,120700,1.5496,1.5496,1.5496,1.5496
20101228,120800,1.5496,1.5496,1.5496,1.5496
20101228,120900,1.5494,1.5494,1.5494,1.5494
20101228,121100,1.5485,1.5485,1.5485,1.5485
20101228,121200,1.5485,1.5485,1.5485,1.5485
20101228,121400,1.5488,1.5488,1.5488,1.5488
20101228,121500,1.5486,1.5486,1.5486,1.5486
20101228,121700,1.5487,1.5487,1.5487,1.5487
20101228,121800,1.5485,1.5485,1.5485,1.5485
20101228,122000,1.5487,1.5487,1.5487,1.5487
20101228,122200,1.5485,1.5485,1.5485,1.5485
20101228,122400,1.5484,1.5484,1.5484,1.5484
20101228,122500,1.5484,1.5484,1.5483,1.5483
20101228,122600,1.5483,1.5483,1.5483,1.5483
20101228,122800,1.5484,1.5486,1.5484,1.5486
20101228,122900,1.5486,1.5486,1.5486,1.5486
20101228,123000,1.5488,1.5488,1.5488,1.5488
20101228,123100,1.5487,1.5487,1.5487,1.5487
20101228,123200,1.5483,1.5483,1.5483,1.5483
20101228,123400,1.5479,1.5479,1.5479,1.5479
20101228,123500,1.548,1.548,1.548,1.548
20101228,123600,1.5482,1.5482,1.5482,1.5482
20101228,123800,1.5482,1.5482,1.5482,1.5482
20101228,123900,1.548,1.548,1.548,1.548
20101228,124000,1.5479,1.5479,1.5479,1.5479
20101228,124100,1.5482,1.5482,1.5482,1.5482
20101228,124300,1.5481,1.5483,1.5481,1.5483
20101228,124400,1.5482,1.5482,1.5482,1.5482
20101228,124500,1.5483,1.5483,1.5483,1.5483
20101228,124600,1.5484,1.5484,1.5484,1.5484
20101228,124800,1.5481,1.5481,1.5481,1.5481
20101228,125000,1.548,1.548,1.5479,1.5479
20101228,125100,1.548,1.548,1.548,1.548
20101228,125200,1.5478,1.5478,1.5478,1.5478
20101228,125300,1.5475,1.5475,1.5475,1.5475
20101228,125400,1.5478,1.5478,1.5478,1.5478
20101228,125500,1.5475,1.5475,1.5475,1.5475
20101228,125600,1.5471,1.5471,1.5471,1.5471
20101228,125800,1.5469,1.5469,1.5469,1.5469
20101228,125900,1.547,1.547,1.547,1.547
20101228,130000,1.547,1.547,1.547,1.547
20101228,130100,1.547,1.547,1.547,1.547
20101228,130200,1.5471,1.5471,1.5471,1.5471
20101228,130400,1.5469,1.5469,1.5469,1.5469
20101228,130500,1.547,1.547,1.547,1.547
20101228,130600,1.547,1.547,1.547,1.547
20101228,130800,1.547,1.5471,1.547,1.5471
20101228,130900,1.5468,1.5468,1.5468,1.5468
20101228,131100,1.5462,1.5462,1.5462,1.5462
20101228,131300,1.5468,1.5468,1.5468,1.5468
20101228,131500,1.5458,1.5458,1.5458,1.5458
20101228,131700,1.546,1.546,1.546,1.546
20101228,131800,1.5464,1.5464,1.5464,1.5464
20101228,131900,1.5461,1.5461,1.5461,1.5461
20101228,132000,1.5464,1.5464,1.5464,1.5464
20101228,132200,1.5468,1.5468,1.5468,1.5468
20101228,132300,1.5475,1.5475,1.5475,1.5475
20101228,132400,1.548,1.548,1.548,1.548
20101228,132500,1.5481,1.5481,1.5481,1.5481
20101228,132700,1.5482,1.5482,1.5482,1.5482
20101228,132800,1.5478,1.5478,1.5478,1.5478
20101228,132900,1.5483,1.5483,1.5483,1.5483
20101228,133000,1.5483,1.5483,1.5483,1.5483
20101228,133100,1.5482,1.5482,1.5482,1.5482
20101228,133300,1.5478,1.5478,1.5478,1.5478
20101228,133400,1.5477,1.5477,1.5477,1.5477
20101228,133500,1.548,1.548,1.548,1.548
20101228,133600,1.5481,1.5481,1.5481,1.5481
20101228,133800,1.5483,1.5483,1.5483,1.5483
20101228,133900,1.5483,1.5483,1.5483,1.5483
20101228,134000,1.5483,1.5483,1.5483,1.5483
20101228,134100,1.5482,1.5482,1.5482,1.5482
20101228,134200,1.5479,1.5479,1.5479,1.5479
20101228,134300,1.5479,1.5479,1.5479,1.5479
20101228,134400,1.5479,1.5479,1.5479,1.5479
20101228,134600,1.5481,1.5481,1.5481,1.5481
20101228,134700,1.548,1.548,1.548,1.548
20101228,134900,1.5476,1.5476,1.5476,1.5476
20101228,135000,1.5476,1.5476,1.5476,1.5476
20101228,135200,1.547,1.547,1.547,1.547
20101228,135300,1.5472,1.5472,1.5472,1.5472
20101228,135500,1.5472,1.5472,1.5472,1.5472
20101228,135600,1.5472,1.5472,1.5472,1.5472
20101228,135800,1.5472,1.5472,1.5471,1.5472
20101228,135900,1.5472,1.5473,1.5472,1.5473
20101228,140000,1.5472,1.5472,1.5472,1.5472
20101228,140100,1.5474,1.5474,1.5474,1.5474
20101228,140200,1.5474,1.5474,1.5474,1.5474
20101228,140300,1.5477,1.5477,1.5477,1.5477
20101228,140400,1.5474,1.5474,1.5474,1.5474
20101228,140600,1.5464,1.5464,1.5464,1.5464
20101228,140800,1.5463,1.5463,1.5463,1.5463
20101228,140900,1.5458,1.5458,1.5458,1.5458
20101228,141100,1.5457,1.5457,1.5457,1.5457
20101228,141200,1.5448,1.5448,1.5448,1.5448
20101228,141400,1.545,1.545,1.545,1.545
20101228,141500,1.5448,1.5448,1.5448,1.5448
20101228,141700,1.5446,1.5446,1.5435,1.5435
20101228,141800,1.5439,1.5439,1.5439,1.5439
20101228,142000,1.5438,1.5443,1.5438,1.5443
20101228,142100,1.5442,1.5442,1.5441,1.5442
20101228,142200,1.5439,1.5439,1.5439,1.5439
20101228,142400,1.544,1.5441,1.5438,1.5438
20101228,142500,1.5434,1.5434,1.5434,1.5434
20101228,142600,1.5432,1.5432,1.5432,1.5432
20101228,142700,1.5431,1.5431,1.5431,1.5431
20101228,142800,1.5426,1.5426,1.5426,1.5426
20101228,142900,1.5417,1.5417,1.5417,1.5417
20101228,143000,1.541,1.541,1.541,1.541
20101228,143100,1.5413,1.5413,1.5413,1.5413
20101228,143200,1.5414,1.5414,1.5414,1.5414
20101228,143300,1.5388,1.5388,1.5388,1.5388
20101228,143400,1.5391,1.5391,1.5391,1.5391
20101228,143500,1.5392,1.5392,1.5392,1.5392
20101228,143600,1.5393,1.5393,1.5393,1.5393
20101228,143800,1.5386,1.5386,1.5386,1.5386
20101228,143900,1.5385,1.5385,1.5385,1.5385
20101228,144000,1.5381,1.5381,1.5381,1.5381
20101228,144100,1.5387,1.5387,1.5387,1.5387
20101228,144200,1.5397,1.5397,1.5397,1.5397
20101228,144300,1.5396,1.5396,1.5396,1.5396
20101228,144400,1.5389,1.5389,1.5389,1.5389
20101228,144500,1.5385,1.5385,1.5385,1.5385
20101228,144600,1.5385,1.5385,1.5385,1.5385
20101228,144700,1.5384,1.5384,1.5384,1.5384
20101228,144800,1.5383,1.5383,1.5383,1.5383
20101228,144900,1.5384,1.5384,1.5384,1.5384
20101228,145000,1.5386,1.5386,1.5386,1.5386
20101228,145100,1.5386,1.5386,1.5386,1.5386
20101228,145200,1.5384,1.5384,1.5384,1.5384
20101228,145300,1.538,1.538,1.538,1.538
20101228,145400,1.538,1.538,1.538,1.538
20101228,145500,1.538,1.538,1.538,1.538
20101228,145600,1.5381,1.5381,1.5381,1.5381
20101228,145800,1.5385,1.5385,1.5385,1.5385
20101228,145900,1.5381,1.5381,1.5381,1.5381
20101228,150000,1.5384,1.5384,1.5384,1.5384
20101228,150100,1.5389,1.5389,1.5389,1.5389
20101228,150200,1.539,1.539,1.539,1.539
20101228,150300,1.5386,1.5386,1.5386,1.5386
20101228,150400,1.5386,1.5386,1.5386,1.5386
20101228,150600,1.5373,1.5373,1.5373,1.5373
20101228,150700,1.5369,1.5369,1.5369,1.5369
20101228,150900,1.5371,1.5371,1.5371,1.5371
20101228,151000,1.5376,1.5376,1.5376,1.5376
20101228,151100,1.5379,1.5379,1.5379,1.5379
20101228,151200,1.538,1.538,1.538,1.538
20101228,151300,1.5379,1.5379,1.5379,1.5379
20101228,151400,1.5376,1.5376,1.5376,1.5376
20101228,151500,1.5374,1.5374,1.5374,1.5374
20101228,151600,1.5374,1.5374,1.5374,1.5374
20101228,151700,1.5378,1.5378,1.5378,1.5378
20101228,151800,1.5377,1.5377,1.5377,1.5377
20101228,151900,1.5385,1.5385,1.5385,1.5385
20101228,152000,1.5384,1.5384,1.5384,1.5384
20101228,152100,1.538,1.538,1.538,1.538
20101228,152200,1.538,1.538,1.538,1.538
20101228,152300,1.5383,1.5383,1.5383,1.5383
20101228,152500,1.5382,1.5384,1.538,1.5384
20101228,152600,1.5383,1.5383,1.5383,1.5383
20101228,152800,1.5384,1.5384,1.5382,1.5383
20101228,152900,1.5386,1.5386,1.5386,1.5386
20101228,153100,1.5387,1.5387,1.5387,1.5387
20101228,153200,1.5385,1.5385,1.5385,1.5385
20101228,153300,1.5386,1.5386,1.5386,1.5386
20101228,153500,1.5385,1.5386,1.5385,1.5385
20101228,153600,1.5386,1.5386,1.5386,1.5386
20101228,153700,1.5385,1.5385,1.5385,1.5385
20101228,153800,1.5385,1.5385,1.5385,1.5385
20101228,154000,1.5387,1.5387,1.5387,1.5387
20101228,154200,1.5386,1.5387,1.5386,1.5386
20101228,154300,1.5389,1.5389,1.5389,1.5389
20101228,154400,1.5387,1.5387,1.5387,1.5387
20101228,154600,1.5388,1.5389,1.5388,1.5388
20101228,154700,1.5391,1.5391,1.5391,1.5391
20101228,154800,1.5391,1.5391,1.5391,1.5391
20101228,154900,1.5389,1.5389,1.5389,1.5389
20101228,155000,1.539,1.539,1.539,1.539
20101228,155200,1.5389,1.5389,1.5387,1.5387
20101228,155300,1.5384,1.5384,1.5384,1.5384
20101228,155400,1.5384,1.5384,1.5384,1.5384
20101228,155500,1.5384,1.5384,1.5384,1.5384
20101228,155600,1.5382,1.5382,1.5382,1.5382
20101228,155800,1.5379,1.5379,1.5379,1.5379
20101228,160000,1.5374,1.5374,1.5374,1.5374
20101228,160200,1.5373,1.5374,1.5372,1.5374
20101228,160300,1.5373,1.5373,1.5369,1.5369
20101228,160400,1.537,1.537,1.537,1.537
20101228,160500,1.5361,1.5361,1.5361,1.5361
20101228,160600,1.536,1.536,1.536,1.536
20101228,160700,1.5359,1.5359,1.5359,1.5359
20101228,160800,1.5359,1.5359,1.5359,1.5359
20101228,161000,1.5361,1.5361,1.5361,1.5361
20101228,161200,1.5365,1.5365,1.5365,1.5365
20101228,161300,1.536,1.536,1.536,1.536
20101228,161500,1.5366,1.5366,1.5366,1.5366
20101228,161600,1.5368,1.5368,1.5368,1.5368
20101228,161700,1.5365,1.5365,1.5365,1.5365
20101228,161800,1.5364,1.5364,1.5364,1.5364
20101228,162000,1.5363,1.5365,1.5362,1.5365
20101228,162100,1.536,1.536,1.536,1.536
20101228,162200,1.536,1.536,1.536,1.536
20101228,162300,1.5363,1.5363,1.5363,1.5363
20101228,162500,1.5364,1.5364,1.5363,1.5364
20101228,162600,1.5359,1.5359,1.5359,1.5359
20101228,162700,1.536,1.536,1.536,1.536
20101228,162800,1.5357,1.5357,1.5357,1.5357
20101228,162900,1.5357,1.5357,1.5357,1.5357
20101228,163000,1.5357,1.5357,1.5357,1.5357
20101228,163200,1.5343,1.5343,1.5343,1.5343
20101228,163300,1.5352,1.5352,1.5352,1.5352
20101228,163500,1.5352,1.5352,1.5349,1.5349
20101228,163600,1.5354,1.5354,1.5354,1.5354
20101228,163700,1.5353,1.5353,1.5353,1.5353
20101228,163900,1.5355,1.5355,1.5355,1.5355
20101228,164000,1.5358,1.5358,1.5358,1.5358
20101228,164100,1.5358,1.5358,1.5358,1.5358
20101228,164200,1.5361,1.5361,1.5361,1.5361
20101228,164300,1.5362,1.5362,1.5362,1.5362
20101228,164400,1.5364,1.5364,1.5364,1.5364
20101228,164500,1.5363,1.5363,1.5363,1.5363
20101228,164700,1.5356,1.5356,1.5356,1.5356
20101228,164800,1.5356,1.5356,1.5356,1.5356
20101228,165000,1.5355,1.5355,1.5354,1.5354
20101228,165100,1.5359,1.5359,1.5359,1.5359
20101228,165200,1.5361,1.5361,1.5361,1.5361
20101228,165400,1.5364,1.5364,1.5364,1.5364
20101228,165500,1.5364,1.5364,1.5364,1.5364
20101228,165700,1.5364,1.5365,1.5364,1.5365
20101228,165800,1.5365,1.5366,1.5365,1.5365
20101228,165900,1.5357,1.5357,1.5357,1.5357
20101228,170100,1.5357,1.5357,1.5357,1.5357
20101228,170300,1.5356,1.5356,1.5356,1.5356
20101228,170500,1.5356,1.5357,1.5355,1.5355
20101228,170600,1.5356,1.5356,1.5356,1.5356
20101228,170700,1.5361,1.5361,1.5361,1.5361
20101228,170900,1.5361,1.5361,1.536,1.536
20101228,171000,1.5359,1.5359,1.5358,1.5358
20101228,171100,1.5362,1.5362,1.5362,1.5362
20101228,171300,1.5361,1.5361,1.536,1.536
20101228,171400,1.5359,1.5362,1.5359,1.5362
20101228,171500,1.536,1.536,1.536,1.536
20101228,171600,1.5359,1.5359,1.5359,1.5359
20101228,171700,1.5356,1.5356,1.5356,1.5356
20101228,171800,1.5366,1.5366,1.5366,1.5366
20101228,172000,1.5365,1.5366,1.5365,1.5366
20101228,172100,1.5372,1.5372,1.5372,1.5372
20101228,172200,1.5373,1.5373,1.5373,1.5373
20101228,172400,1.5372,1.5372,1.5372,1.5372
20101228,172500,1.5373,1.5374,1.5372,1.5374
20101228,172600,1.5375,1.5375,1.5375,1.5375
20101228,172700,1.5377,1.5377,1.5377,1.5377
20101228,172800,1.5384,1.5384,1.5384,1.5384
20101228,172900,1.5384,1.5384,1.5384,1.5384
20101228,173000,1.5385,1.5385,1.5385,1.5385
20101228,173100,1.5384,1.5384,1.5384,1.5384
20101228,173300,1.5388,1.5388,1.5388,1.5388
20101228,173500,1.5386,1.5386,1.5386,1.5386
20101228,173700,1.5386,1.5386,1.5385,1.5386
20101228,173800,1.5387,1.5387,1.5384,1.5384
20101228,173900,1.5383,1.5383,1.5383,1.5383
20101228,174000,1.5384,1.5384,1.5384,1.5384
20101228,174100,1.5384,1.5384,1.5384,1.5384
20101228,174200,1.5383,1.5383,1.5383,1.5383
20101228,174400,1.5383,1.5384,1.5383,1.5383
20101228,174500,1.5383,1.5384,1.5383,1.5383
20101228,174600,1.5382,1.5382,1.5382,1.5382
20101228,174800,1.5381,1.5381,1.5381,1.5381
20101228,175000,1.538,1.538,1.538,1.538
20101228,175100,1.5381,1.5381,1.5381,1.5381
20101228,175300,1.5379,1.5379,1.5379,1.5379
20101228,175400,1.5379,1.5379,1.5379,1.5379
20101228,175600,1.5379,1.5379,1.5379,1.5379
20101228,175700,1.5378,1.5378,1.5378,1.5378
20101228,175800,1.5377,1.5377,1.5377,1.5377
20101228,180000,1.5378,1.5379,1.5377,1.5379
20101228,180100,1.538,1.538,1.5379,1.5379
20101228,180200,1.5379,1.5379,1.5372,1.5372
20101228,180300,1.5373,1.5373,1.5369,1.5369
20101228,180400,1.5368,1.5368,1.5365,1.5368
20101228,180500,1.5368,1.5368,1.5365,1.5365
20101228,180600,1.5364,1.5364,1.5364,1.5364
20101228,180700,1.5365,1.5365,1.5364,1.5365
20101228,180800,1.5365,1.5365,1.5365,1.5365
20101228,180900,1.5365,1.5369,1.5365,1.5369
20101228,181000,1.5369,1.5369,1.5368,1.5368
20101228,181100,1.5367,1.5367,1.5364,1.5365
20101228,181200,1.5365,1.5365,1.5364,1.5365
20101228,181300,1.5365,1.5365,1.5363,1.5364
20101228,181400,1.5364,1.5368,1.5364,1.5368
20101228,181500,1.5367,1.5371,1.5367,1.537
20101228,181600,1.5371,1.5371,1.5368,1.537
20101228,181700,1.5371,1.5371,1.537,1.537
20101228,181800,1.537,1.537,1.5367,1.5367
20101228,181900,1.5366,1.5366,1.5365,1.5366
20101228,182000,1.5365,1.5365,1.5365,1.5365
20101228,182100,1.5364,1.5364,1.5363,1.5363
20101228,182200,1.5362,1.5362,1.536,1.536
20101228,182300,1.536,1.5361,1.536,1.5361
20101228,182400,1.536,1.536,1.536,1.536
20101228,182500,1.536,1.5361,1.5359,1.5361
20101228,182600,1.536,1.5361,1.536,1.536
20101228,182700,1.5361,1.5361,1.536,1.5361
20101228,182800,1.5362,1.5362,1.5361,1.5361
20101228,182900,1.5361,1.5361,1.536,1.5361
20101228,183000,1.536,1.5361,1.5359,1.536
20101228,183100,1.5361,1.5361,1.536,1.5361
20101228,183200,1.5361,1.5361,1.5361,1.5361
20101228,183300,1.5361,1.5361,1.536,1.536
20101228,183400,1.5361,1.5364,1.5361,1.5364
20101228,183500,1.5363,1.5363,1.5359,1.5359
20101228,183600,1.5358,1.5358,1.5356,1.5357
20101228,183700,1.5358,1.5359,1.5358,1.5359
20101228,183800,1.536,1.5361,1.5359,1.5359
20101228,183900,1.536,1.536,1.5358,1.5359
20101228,184000,1.536,1.5361,1.536,1.536
20101228,184100,1.536,1.536,1.5357,1.5358
20101228,184200,1.5357,1.5358,1.5357,1.5357
20101228,184300,1.5357,1.5358,1.5357,1.5357
20101228,184400,1.5357,1.5359,1.5357,1.5359
20101228,184500,1.5358,1.5358,1.5357,1.5357
20101228,184600,1.5358,1.5358,1.5356,1.5356
20101228,184700,1.5356,1.5356,1.5356,1.5356
20101228,184800,1.5355,1.5356,1.5355,1.5355
20101228,184900,1.5354,1.5355,1.5353,1.5353
20101228,185000,1.5353,1.5353,1.5352,1.5353
20101228,185100,1.5353,1.5353,1.5352,1.5353
20101228,185200,1.5354,1.5355,1.5354,1.5355
20101228,185300,1.5354,1.5355,1.5354,1.5354
20101228,185400,1.5354,1.5354,1.5353,1.5353
20101228,185500,1.5353,1.5353,1.5353,1.5353
20101228,185600,1.5353,1.5353,1.5353,1.5353
20101228,185700,1.5352,1.5354,1.5352,1.5353
20101228,185800,1.5353,1.5353,1.5353,1.5353
20101228,185900,1.5353,1.5353,1.5353,1.5353
20101228,190000,1.5352,1.5353,1.5352,1.5353
20101228,190100,1.5353,1.5353,1.5352,1.5352
20101228,190200,1.5352,1.5353,1.5352,1.5353
20101228,190300,1.5354,1.5357,1.5353,1.5356
20101228,190400,1.5356,1.5358,1.5355,1.5358
20101228,190500,1.5357,1.5358,1.5357,1.5358
20101228,190600,1.5358,1.536,1.5358,1.536
20101228,190700,1.5361,1.5362,1.5361,1.5362
20101228,190800,1.5363,1.5365,1.5363,1.5365
20101228,190900,1.5364,1.5367,1.5364,1.5367
20101228,191000,1.5368,1.5368,1.5365,1.5365
20101228,191100,1.5366,1.5368,1.5366,1.5368
20101228,191200,1.5369,1.5371,1.5368,1.5371
20101228,191300,1.5372,1.5374,1.537,1.5374
20101228,191400,1.5375,1.5377,1.5375,1.5376
20101228,191500,1.5377,1.5377,1.5373,1.5373
20101228,191600,1.5374,1.5375,1.5374,1.5375
20101228,191700,1.5376,1.5376,1.5375,1.5375
20101228,191800,1.5376,1.5376,1.5375,1.5375
20101228,191900,1.5375,1.5375,1.5374,1.5374
20101228,192000,1.5374,1.5374,1.5372,1.5372
20101228,192100,1.5372,1.5374,1.5372,1.5374
20101228,192200,1.5374,1.5375,1.5374,1.5374
20101228,192300,1.5375,1.5376,1.5375,1.5376
20101228,192400,1.5376,1.5377,1.5376,1.5376
20101228,192500,1.5376,1.5376,1.5376,1.5376
20101228,192600,1.5376,1.5377,1.5376,1.5377
20101228,192700,1.5376,1.5377,1.5375,1.5375
20101228,192800,1.5375,1.5375,1.5375,1.5375
20101228,192900,1.5375,1.5376,1.5375,1.5376
20101228,193000,1.5375,1.5375,1.5374,1.5374
20101228,193100,1.5374,1.5374,1.5373,1.5373
20101228,193200,1.5373,1.5373,1.5372,1.5372
20101228,193300,1.5372,1.5373,1.5372,1.5373
20101228,193400,1.5374,1.5374,1.5373,1.5374
20101228,193500,1.5374,1.5376,1.5374,1.5376
20101228,193600,1.5376,1.5376,1.5375,1.5376
20101228,193700,1.5375,1.5376,1.5375,1.5376
20101228,193800,1.5375,1.5376,1.5375,1.5375
20101228,193900,1.5375,1.5375,1.5374,1.5374
20101228,194000,1.5373,1.5374,1.5373,1.5374
20101228,194100,1.5374,1.5374,1.5374,1.5374
20101228,194200,1.5373,1.5374,1.5372,1.5373
20101228,194300,1.5372,1.5372,1.5372,1.5372
20101228,194400,1.5372,1.5373,1.5372,1.5372
20101228,194500,1.5371,1.5371,1.537,1.537
20101228,194600,1.537,1.5371,1.537,1.5371
20101228,194700,1.5371,1.5371,1.5371,1.5371
20101228,194800,1.5371,1.5371,1.5371,1.5371
20101228,194900,1.5371,1.5371,1.537,1.537
20101228,195000,1.537,1.5371,1.537,1.5371
20101228,195100,1.5372,1.5372,1.5371,1.5372
20101228,195200,1.5372,1.5372,1.5372,1.5372
20101228,195300,1.5371,1.5372,1.537,1.537
20101228,195400,1.5369,1.5369,1.5367,1.5368
20101228,195500,1.5369,1.5371,1.5369,1.5371
20101228,195600,1.5371,1.5372,1.537,1.537
20101228,195700,1.5371,1.5371,1.5369,1.5369
20101228,195800,1.537,1.5372,1.537,1.5372
20101228,195900,1.5373,1.5373,1.5372,1.5372
20101228,200000,1.5371,1.5371,1.5368,1.5368
20101228,200100,1.5369,1.5371,1.5369,1.5371
20101228,200200,1.5372,1.5372,1.5372,1.5372
20101228,200300,1.5372,1.5372,1.5371,1.5371
20101228,200400,1.5372,1.5372,1.5371,1.5371
20101228,200500,1.5371,1.5371,1.5371,1.5371
20101228,200600,1.5372,1.5373,1.5371,1.5372
20101228,200700,1.5372,1.5372,1.5371,1.5371
20101228,200800,1.5372,1.5373,1.5372,1.5372
20101228,200900,1.5371,1.5371,1.5371,1.5371
20101228,201000,1.537,1.5371,1.537,1.5371
20101228,201100,1.537,1.5371,1.537,1.537
20101228,201200,1.537,1.5371,1.537,1.5371
20101228,201300,1.5371,1.5371,1.5371,1.5371
20101228,201400,1.5371,1.5372,1.5371,1.5372
20101228,201500,1.5371,1.5372,1.5371,1.5372
20101228,201600,1.5372,1.5373,1.5372,1.5372
20101228,201700,1.5372,1.5372,1.5372,1.5372
20101228,201800,1.5372,1.5372,1.5371,1.5372
20101228,201900,1.5371,1.5371,1.5371,1.5371
20101228,202000,1.5371,1.5371,1.537,1.537
20101228,202100,1.5371,1.5371,1.5369,1.5369
20101228,202200,1.537,1.5371,1.537,1.537
20101228,202300,1.537,1.537,1.537,1.537
20101228,202400,1.537,1.537,1.537,1.537
20101228,202500,1.537,1.537,1.537,1.537
20101228,202600,1.537,1.5371,1.537,1.537
20101228,202700,1.537,1.5371,1.537,1.5371
20101228,202800,1.5371,1.5371,1.5371,1.5371
20101228,202900,1.5371,1.5371,1.5371,1.5371
20101228,203000,1.5371,1.5372,1.5371,1.5372
20101228,203100,1.5372,1.5372,1.5372,1.5372
20101228,203200,1.5371,1.5372,1.5371,1.5372
20101228,203300,1.5373,1.5374,1.5373,1.5374
20101228,203400,1.5374,1.5374,1.5373,1.5374
20101228,203500,1.5374,1.5374,1.5372,1.5373
20101228,203600,1.5372,1.5373,1.5372,1.5372
20101228,203700,1.5372,1.5373,1.5372,1.5372
20101228,203800,1.5373,1.5374,1.5372,1.5374
20101228,203900,1.5375,1.5377,1.5375,1.5377
20101228,204000,1.5376,1.5376,1.5376,1.5376
20101228,204100,1.5376,1.5376,1.5376,1.5376
20101228,204200,1.5376,1.5377,1.5376,1.5376
20101228,204300,1.5377,1.5377,1.5377,1.5377
20101228,204400,1.5377,1.5379,1.5377,1.5379
20101228,204500,1.5379,1.538,1.5379,1.5379
20101228,204600,1.538,1.5381,1.5379,1.5381
20101228,204700,1.538,1.5381,1.538,1.538
20101228,204800,1.5381,1.5381,1.538,1.5381
20101228,204900,1.5381,1.5381,1.5381,1.5381
20101228,205000,1.5381,1.5381,1.5381,1.5381
20101228,205100,1.5382,1.5382,1.5381,1.5381
20101228,205200,1.5381,1.5381,1.5381,1.5381
20101228,205300,1.538,1.5381,1.538,1.538
20101228,205400,1.538,1.538,1.538,1.538
20101228,205500,1.5379,1.5381,1.5379,1.5381
20101228,205600,1.5382,1.5382,1.5381,1.5381
20101228,205700,1.5382,1.5383,1.5382,1.5383
20101228,205800,1.5383,1.5383,1.5383,1.5383
20101228,205900,1.5383,1.5383,1.5383,1.5383
20101228,210000,1.5383,1.5383,1.5383,1.5383
20101228,210100,1.5383,1.5383,1.5382,1.5382
20101228,210200,1.5383,1.5383,1.5381,1.5381
20101228,210300,1.5381,1.5382,1.538,1.5382
20101228,210400,1.5382,1.5383,1.5382,1.5383
20101228,210500,1.5382,1.5382,1.5382,1.5382
20101228,210600,1.5382,1.5382,1.538,1.538
20101228,210700,1.5379,1.538,1.5379,1.538
20101228,210800,1.538,1.5381,1.538,1.538
20101228,210900,1.538,1.538,1.5379,1.538
20101228,211000,1.538,1.5381,1.538,1.5381
20101228,211100,1.538,1.538,1.538,1.538
20101228,211200,1.538,1.538,1.5378,1.5378
20101228,211300,1.5379,1.538,1.5378,1.538
20101228,211400,1.5381,1.5381,1.5381,1.5381
20101228,211500,1.5381,1.5381,1.5381,1.5381
20101228,211600,1.5381,1.5381,1.5381,1.5381
20101228,211700,1.5381,1.5381,1.5381,1.5381
20101228,211800,1.5381,1.5381,1.5381,1.5381
20101228,211900,1.5382,1.5382,1.5381,1.5381
20101228,212000,1.5381,1.5382,1.5379,1.5379
20101228,212100,1.5379,1.5379,1.5378,1.5378
20101228,212200,1.5378,1.5379,1.5378,1.5378
20101228,212300,1.5378,1.5379,1.5378,1.5378
20101228,212400,1.5378,1.5378,1.5378,1.5378
20101228,212500,1.5378,1.5381,1.5378,1.538
20101228,212600,1.5381,1.5382,1.5381,1.5382
20101228,212700,1.5383,1.5383,1.5382,1.5382
20101228,212800,1.5383,1.5383,1.5382,1.5383
20101228,212900,1.5382,1.5384,1.5382,1.5384
20101228,213000,1.5384,1.5384,1.5384,1.5384
20101228,213100,1.5384,1.5384,1.5383,1.5384
20101228,213200,1.5384,1.5384,1.5384,1.5384
20101228,213300,1.5383,1.5383,1.5382,1.5382
20101228,213400,1.5383,1.5383,1.5382,1.5382
20101228,213500,1.5382,1.5382,1.5381,1.5382
20101228,213600,1.5381,1.5382,1.5381,1.5382
20101228,213700,1.5381,1.5382,1.5381,1.5381
20101228,213800,1.5381,1.5381,1.538,1.5381
20101228,213900,1.5381,1.5381,1.5377,1.5377
20101228,214000,1.5375,1.538,1.5374,1.538
20101228,214100,1.5381,1.5381,1.5381,1.5381
20101228,214200,1.5381,1.5381,1.538,1.5381
20101228,214300,1.538,1.538,1.538,1.538
20101228,214400,1.538,1.538,1.538,1.538
20101228,214500,1.538,1.538,1.5374,1.5374
20101228,214600,1.5375,1.5375,1.5374,1.5374
20101228,214700,1.5374,1.5374,1.5374,1.5374
20101228,214800,1.5373,1.5374,1.5373,1.5374
20101228,214900,1.5374,1.5375,1.5373,1.5374
20101228,215000,1.5373,1.5374,1.5373,1.5374
20101228,215100,1.5374,1.5375,1.5374,1.5374
20101228,215200,1.5373,1.5374,1.5373,1.5374
20101228,215300,1.5373,1.5373,1.5369,1.537
20101228,215400,1.5369,1.537,1.5369,1.5369
20101228,215500,1.5368,1.5368,1.5367,1.5367
20101228,215600,1.5368,1.5368,1.5368,1.5368
20101228,215700,1.5369,1.5371,1.5367,1.5367
20101228,215800,1.5368,1.5369,1.5367,1.5367
20101228,215900,1.5367,1.5367,1.5366,1.5366
20101228,220000,1.5366,1.5366,1.5365,1.5366
20101228,220100,1.5364,1.5365,1.5363,1.5364
20101228,220200,1.5365,1.5366,1.5365,1.5366
20101228,220300,1.5365,1.5365,1.5364,1.5365
20101228,220400,1.5366,1.5369,1.5366,1.5369
20101228,220500,1.5369,1.5369,1.5368,1.5368
20101228,220600,1.5368,1.5368,1.5367,1.5367
20101228,220700,1.5367,1.5368,1.5365,1.5367
20101228,220800,1.5366,1.5369,1.5365,1.5367
20101228,220900,1.5368,1.5369,1.5367,1.5369
20101228,221000,1.5368,1.5368,1.5363,1.5363
20101228,221100,1.5364,1.537,1.5363,1.5369
20101228,221200,1.5368,1.5369,1.5367,1.5369
20101228,221300,1.5369,1.537,1.5366,1.5366
20101228,221400,1.5365,1.5366,1.5365,1.5366
20101228,221500,1.5365,1.5366,1.5364,1.5366
20101228,221600,1.5366,1.5366,1.5365,1.5365
20101228,221700,1.5366,1.5366,1.5364,1.5365
20101228,221800,1.5365,1.5365,1.5365,1.5365
20101228,221900,1.5365,1.5365,1.5364,1.5364
20101228,222000,1.5364,1.5365,1.5364,1.5365
20101228,222100,1.5365,1.5366,1.5365,1.5365
20101228,222200,1.5364,1.5364,1.5362,1.5363
20101228,222300,1.5364,1.5364,1.5363,1.5363
20101228,222400,1.5364,1.5367,1.5364,1.5364
20101228,222500,1.5364,1.5364,1.5364,1.5364
20101228,222600,1.5365,1.5365,1.5363,1.5363
20101228,222700,1.5363,1.5364,1.5363,1.5364
20101228,222800,1.5364,1.5364,1.5364,1.5364
20101228,222900,1.5364,1.5364,1.5363,1.5363
20101228,223000,1.5363,1.5364,1.5363,1.5363
20101228,223100,1.5363,1.5363,1.5362,1.5362
20101228,223200,1.5362,1.5362,1.5361,1.5362
20101228,223300,1.5362,1.5362,1.5361,1.5362
20101228,223400,1.5362,1.5362,1.5362,1.5362
20101228,223500,1.5361,1.5362,1.5361,1.5362
20101228,223600,1.5362,1.5362,1.5362,1.5362
20101228,223700,1.5362,1.5362,1.5362,1.5362
20101228,223800,1.5362,1.5362,1.5362,1.5362
20101228,223900,1.5361,1.5361,1.5357,1.5357
20101228,224000,1.5357,1.5358,1.5357,1.5358
20101228,224100,1.5358,1.5358,1.5357,1.5358
20101228,224200,1.5357,1.5357,1.5357,1.5357
20101228,224400,1.5357,1.5357,1.5357,1.5357
20101228,224500,1.5357,1.5357,1.5357,1.5357
20101228,224600,1.5357,1.5358,1.5357,1.5358
20101228,224700,1.5358,1.5358,1.5358,1.5358
20101228,224900,1.5359,1.5359,1.5359,1.5359
20101228,225100,1.5362,1.5362,1.5362,1.5362
20101228,225200,1.5362,1.5362,1.5362,1.5362
20101228,225400,1.5363,1.5363,1.5362,1.5362
20101228,225500,1.5362,1.5362,1.5362,1.5362
20101228,225600,1.5362,1.5362,1.5362,1.5362
20101228,225800,1.5362,1.5363,1.5362,1.5363
20101228,225900,1.5363,1.5363,1.5363,1.5363
20101228,230000,1.5366,1.5366,1.5366,1.5366
20101228,230100,1.5365,1.5365,1.5365,1.5365
20101228,230200,1.5362,1.5362,1.5362,1.5362
20101228,230400,1.5363,1.5363,1.5363,1.5363
20101228,230500,1.5363,1.5363,1.5363,1.5363
20101228,230600,1.5363,1.5363,1.5363,1.5363
20101228,230700,1.5363,1.5363,1.5363,1.5363
20101228,230900,1.5364,1.5364,1.5363,1.5363
20101228,231000,1.5364,1.5364,1.5363,1.5363
20101228,231100,1.5363,1.5363,1.5363,1.5363
20101228,231200,1.5363,1.5363,1.5363,1.5363
20101228,231300,1.5363,1.5363,1.5363,1.5363
20101228,231400,1.5363,1.5363,1.5363,1.5363
20101228,231600,1.5363,1.5363,1.5363,1.5363
20101228,231700,1.5363,1.5364,1.5363,1.5364
20101228,231800,1.5364,1.5364,1.5364,1.5364
20101228,231900,1.5363,1.5364,1.5363,1.5363
20101228,232000,1.5363,1.5364,1.5363,1.5364
20101228,232100,1.5364,1.5364,1.5363,1.5363
20101228,232200,1.5363,1.5364,1.5363,1.5364
20101228,232300,1.5364,1.5366,1.5364,1.5366
20101228,232400,1.5366,1.5367,1.5366,1.5366
20101228,232500,1.5366,1.5366,1.5366,1.5366
20101228,232700,1.5366,1.5366,1.5366,1.5366
20101228,232900,1.5364,1.5364,1.5364,1.5364
20101228,233100,1.5364,1.5364,1.5364,1.5364
20101228,233300,1.5363,1.5363,1.5363,1.5363
20101228,233500,1.5362,1.5362,1.5362,1.5362
20101228,233600,1.5364,1.5364,1.5364,1.5364
20101228,233800,1.5362,1.5362,1.5362,1.5362
20101228,234000,1.5362,1.5362,1.5362,1.5362
20101228,234100,1.5358,1.5358,1.5358,1.5358
20101228,234200,1.5358,1.5358,1.5358,1.5358
20101228,234300,1.5358,1.5358,1.5358,1.5358
20101228,234400,1.5359,1.5359,1.5359,1.5359
20101228,234500,1.5359,1.5359,1.5359,1.5359
20101228,234700,1.5356,1.5356,1.5356,1.5356
20101228,234800,1.5356,1.5356,1.5356,1.5356
20101228,235000,1.5353,1.5353,1.5353,1.5353
20101228,235100,1.5351,1.5351,1.5351,1.5351
20101228,235200,1.5351,1.5351,1.5351,1.5351
20101228,235400,1.5351,1.5351,1.5351,1.5351
20101228,235600,1.535,1.535,1.535,1.535
20101228,235700,1.5351,1.5351,1.5351,1.5351
20101228,235800,1.5352,1.5352,1.5352,1.5352
20101228,235900,1.5352,1.5352,1.5352,1.5352
20101229,0,1.5352,1.5352,1.5352,1.5352
20101229,100,1.5353,1.5353,1.5353,1.5353
20101229,300,1.5353,1.5356,1.5353,1.5354
20101229,400,1.5355,1.5356,1.5354,1.5354
20101229,500,1.5354,1.5354,1.5352,1.5352
20101229,600,1.5353,1.5354,1.5352,1.5354
20101229,700,1.5353,1.5355,1.5353,1.5354
20101229,800,1.5358,1.5358,1.5358,1.5358
20101229,900,1.5359,1.5359,1.5359,1.5359
20101229,1100,1.536,1.536,1.536,1.536
20101229,1200,1.5361,1.5361,1.5361,1.5361
20101229,1300,1.536,1.536,1.536,1.536
20101229,1500,1.536,1.536,1.536,1.536
20101229,1600,1.5359,1.5359,1.5359,1.5359
20101229,1800,1.536,1.536,1.536,1.536
20101229,1900,1.536,1.536,1.536,1.536
20101229,2100,1.5359,1.5359,1.5359,1.5359
20101229,2300,1.5359,1.536,1.5358,1.536
20101229,2400,1.536,1.536,1.5359,1.5359
20101229,2500,1.5359,1.5359,1.5358,1.5358
20101229,2600,1.5359,1.5359,1.5358,1.5358
20101229,2700,1.5358,1.5359,1.5358,1.5358
20101229,2800,1.5358,1.5359,1.5358,1.5359
20101229,2900,1.5359,1.5359,1.5359,1.5359
20101229,3100,1.5363,1.5363,1.5363,1.5363
20101229,3300,1.5364,1.5372,1.5364,1.5372
20101229,3400,1.5378,1.5378,1.5378,1.5378
20101229,3500,1.5373,1.5373,1.5373,1.5373
20101229,3600,1.5379,1.5379,1.5379,1.5379
20101229,3800,1.5374,1.5374,1.5374,1.5374
20101229,3900,1.5375,1.5375,1.5375,1.5375
20101229,4000,1.538,1.538,1.538,1.538
20101229,4200,1.5384,1.5384,1.5384,1.5384
20101229,4300,1.5387,1.5387,1.5387,1.5387
20101229,4500,1.5386,1.5386,1.5386,1.5386
20101229,4600,1.5386,1.5386,1.5386,1.5386
20101229,4700,1.5385,1.5385,1.5385,1.5385
20101229,4800,1.5383,1.5383,1.5383,1.5383
20101229,5000,1.5384,1.5384,1.5384,1.5384
20101229,5100,1.5384,1.5384,1.5384,1.5384
20101229,5200,1.5385,1.5385,1.5385,1.5385
20101229,5300,1.5383,1.5383,1.5383,1.5383
20101229,5400,1.5383,1.5383,1.5383,1.5383
20101229,5500,1.5384,1.5384,1.5384,1.5384
20101229,5600,1.5383,1.5383,1.5383,1.5383
20101229,5800,1.5382,1.5387,1.5382,1.5383
20101229,5900,1.5384,1.5384,1.5383,1.5383
20101229,10000,1.5382,1.5384,1.5382,1.5383
20101229,10100,1.5383,1.5384,1.5383,1.5384
20101229,10200,1.5383,1.5383,1.5383,1.5383
20101229,10300,1.5383,1.5383,1.5374,1.5376
20101229,10400,1.5384,1.5384,1.5384,1.5384
20101229,10500,1.5383,1.5383,1.5383,1.5383
20101229,10600,1.5383,1.5383,1.5383,1.5383
20101229,10800,1.5388,1.5388,1.5388,1.5388
20101229,11000,1.5389,1.5389,1.5384,1.5387
20101229,11100,1.5387,1.5387,1.5385,1.5385
20101229,11200,1.5384,1.5384,1.5384,1.5384
20101229,11400,1.5383,1.5383,1.5383,1.5383
20101229,11500,1.5384,1.5384,1.5384,1.5384
20101229,11700,1.5384,1.5384,1.5383,1.5383
20101229,11800,1.5383,1.5385,1.5383,1.5385
20101229,11900,1.5384,1.5385,1.5384,1.5384
20101229,12000,1.5383,1.5383,1.5382,1.5382
20101229,12100,1.5382,1.5386,1.5382,1.5386
20101229,12200,1.5385,1.5387,1.5385,1.5385
20101229,12300,1.5384,1.5384,1.5384,1.5384
20101229,12500,1.5386,1.5386,1.5386,1.5386
20101229,12700,1.5388,1.5388,1.5388,1.5388
20101229,12900,1.5388,1.5388,1.5387,1.5387
20101229,13000,1.5388,1.5388,1.5388,1.5388
20101229,13100,1.5388,1.5388,1.5388,1.5388
20101229,13200,1.5388,1.5388,1.5388,1.5388
20101229,13400,1.5388,1.5388,1.5388,1.5388
20101229,13500,1.5388,1.5388,1.5388,1.5388
20101229,13600,1.5389,1.5389,1.5389,1.5389
20101229,13700,1.5385,1.5385,1.5385,1.5385
20101229,13900,1.5385,1.5385,1.5385,1.5385
20101229,14000,1.5384,1.5384,1.5384,1.5384
20101229,14100,1.5384,1.5384,1.5384,1.5384
20101229,14200,1.5384,1.5384,1.5384,1.5384
20101229,14400,1.5384,1.5384,1.5383,1.5383
20101229,14500,1.5384,1.5384,1.5384,1.5384
20101229,14700,1.5384,1.5384,1.5384,1.5384
20101229,14800,1.5384,1.5384,1.5384,1.5384
20101229,14900,1.5384,1.5384,1.5384,1.5384
20101229,15000,1.5383,1.5383,1.5383,1.5383
20101229,15100,1.5383,1.5383,1.5383,1.5383
20101229,15200,1.5386,1.5386,1.5386,1.5386
20101229,15400,1.5387,1.5387,1.5387,1.5387
20101229,15500,1.5389,1.5389,1.5389,1.5389
20101229,15600,1.539,1.539,1.539,1.539
20101229,15700,1.5389,1.5389,1.5389,1.5389
20101229,15800,1.539,1.539,1.539,1.539
20101229,15900,1.539,1.539,1.539,1.539
20101229,20000,1.5391,1.5391,1.5391,1.5391
20101229,20100,1.5391,1.5391,1.5391,1.5391
20101229,20200,1.5392,1.5392,1.5392,1.5392
20101229,20400,1.5389,1.5389,1.5389,1.5389
20101229,20600,1.539,1.539,1.5389,1.539
20101229,20700,1.5391,1.5391,1.5391,1.5391
20101229,20800,1.5391,1.5392,1.5391,1.5391
20101229,20900,1.5392,1.5392,1.539,1.539
20101229,21000,1.5391,1.5391,1.5391,1.5391
20101229,21100,1.5391,1.5391,1.5391,1.5391
20101229,21200,1.5391,1.5391,1.5391,1.5391
20101229,21300,1.5391,1.5391,1.5391,1.5391
20101229,21500,1.5391,1.5391,1.5391,1.5391
20101229,21600,1.5391,1.5391,1.539,1.539
20101229,21700,1.539,1.539,1.539,1.539
20101229,21900,1.539,1.539,1.539,1.539
20101229,22100,1.5391,1.5391,1.5391,1.5391
20101229,22200,1.5392,1.5392,1.5392,1.5392
20101229,22300,1.5393,1.5393,1.5393,1.5393
20101229,22500,1.5392,1.5392,1.5392,1.5392
20101229,22700,1.5392,1.5392,1.5391,1.5392
20101229,22800,1.5394,1.5394,1.5394,1.5394
20101229,22900,1.5394,1.5394,1.5394,1.5394
20101229,23000,1.5393,1.5393,1.5393,1.5393
20101229,23100,1.5393,1.5393,1.5393,1.5393
20101229,23200,1.5395,1.5395,1.5395,1.5395
20101229,23300,1.5396,1.5396,1.5396,1.5396
20101229,23500,1.5395,1.5398,1.5395,1.5398
20101229,23600,1.5399,1.5399,1.5399,1.5399
20101229,23800,1.54,1.54,1.5398,1.5399
20101229,23900,1.5399,1.54,1.5399,1.54
20101229,24000,1.54,1.54,1.5399,1.5399
20101229,24100,1.5399,1.5399,1.5399,1.5399
20101229,24200,1.5397,1.5397,1.5397,1.5397
20101229,24400,1.5398,1.5398,1.5398,1.5398
20101229,24600,1.5398,1.5398,1.5398,1.5398
20101229,24700,1.5397,1.5398,1.5397,1.5398
20101229,24800,1.5398,1.5398,1.5397,1.5397
20101229,24900,1.5397,1.5398,1.5397,1.5397
20101229,25000,1.5397,1.5397,1.5397,1.5397
20101229,25100,1.5395,1.5395,1.5395,1.5395
20101229,25300,1.5394,1.5394,1.5394,1.5394
20101229,25400,1.5392,1.5392,1.5392,1.5392
20101229,25500,1.5392,1.5392,1.5392,1.5392
20101229,25700,1.5393,1.5393,1.5393,1.5393
20101229,25800,1.5394,1.5394,1.5394,1.5394
20101229,25900,1.5396,1.5396,1.5396,1.5396
20101229,30000,1.5399,1.5399,1.5399,1.5399
20101229,30200,1.5399,1.5399,1.5399,1.5399
20101229,30400,1.5399,1.54,1.5399,1.54
20101229,30500,1.5398,1.5398,1.5398,1.5398
20101229,30600,1.5397,1.5397,1.5397,1.5397
20101229,30800,1.5398,1.5398,1.5397,1.5398
20101229,30900,1.5398,1.5398,1.5398,1.5398
20101229,31000,1.5398,1.5399,1.5398,1.5399
20101229,31100,1.54,1.54,1.5399,1.5399
20101229,31200,1.54,1.54,1.5399,1.5399
20101229,31300,1.5399,1.5399,1.5399,1.5399
20101229,31500,1.5401,1.5401,1.5401,1.5401
20101229,31600,1.5401,1.5401,1.5401,1.5401
20101229,31700,1.5402,1.5402,1.5402,1.5402
20101229,31800,1.5402,1.5402,1.5402,1.5402
20101229,31900,1.5402,1.5402,1.5402,1.5402
20101229,32000,1.5401,1.5401,1.5401,1.5401
20101229,32200,1.5401,1.5401,1.54,1.54
20101229,32300,1.54,1.54,1.54,1.54
20101229,32400,1.54,1.54,1.54,1.54
20101229,32500,1.54,1.54,1.54,1.54
20101229,32600,1.5399,1.5399,1.5398,1.5398
20101229,32700,1.5398,1.5398,1.5396,1.5396
20101229,32800,1.5397,1.5397,1.5388,1.5394
20101229,32900,1.5393,1.5396,1.5393,1.5395
20101229,33000,1.5393,1.5393,1.5393,1.5393
20101229,33200,1.5393,1.5393,1.5393,1.5393
20101229,33400,1.5393,1.5393,1.5393,1.5393
20101229,33500,1.5393,1.5393,1.5393,1.5393
20101229,33600,1.5393,1.5393,1.5393,1.5393
20101229,33700,1.5393,1.5393,1.5393,1.5393
20101229,33800,1.5392,1.5392,1.5392,1.5392
20101229,33900,1.5393,1.5393,1.5393,1.5393
20101229,34000,1.5394,1.5394,1.5394,1.5394
20101229,34100,1.5395,1.5395,1.5395,1.5395
20101229,34300,1.5393,1.5393,1.5393,1.5393
20101229,34500,1.5392,1.5393,1.5392,1.5393
20101229,34600,1.5395,1.5395,1.5395,1.5395
20101229,34800,1.5395,1.5395,1.5394,1.5394
20101229,34900,1.5395,1.5395,1.5395,1.5395
20101229,35000,1.5395,1.5395,1.5393,1.5393
20101229,35100,1.5393,1.5393,1.5393,1.5393
20101229,35200,1.5394,1.5394,1.5394,1.5394
20101229,35300,1.5393,1.5393,1.5393,1.5393
20101229,35400,1.5394,1.5394,1.5394,1.5394
20101229,35600,1.5394,1.5394,1.5393,1.5393
20101229,35700,1.5393,1.5396,1.5393,1.5396
20101229,35800,1.5396,1.5396,1.5394,1.5394
20101229,35900,1.5395,1.5395,1.5395,1.5395
20101229,40100,1.5395,1.5395,1.5394,1.5395
20101229,40200,1.5395,1.5397,1.5395,1.5395
20101229,40300,1.5396,1.5397,1.5396,1.5397
20101229,40400,1.5398,1.5398,1.5398,1.5398
20101229,40600,1.5398,1.5398,1.5398,1.5398
20101229,40700,1.54,1.54,1.54,1.54
20101229,40900,1.54,1.5401,1.54,1.54
20101229,41000,1.54,1.54,1.54,1.54
20101229,41100,1.54,1.54,1.54,1.54
20101229,41200,1.5399,1.5399,1.5399,1.5399
20101229,41400,1.5398,1.5401,1.5398,1.5401
20101229,41500,1.5401,1.5401,1.54,1.5401
20101229,41600,1.5401,1.5401,1.54,1.54
20101229,41700,1.5401,1.5401,1.5401,1.5401
20101229,41800,1.5401,1.5401,1.5401,1.5401
20101229,41900,1.5403,1.5403,1.5403,1.5403
20101229,42000,1.5403,1.5403,1.5403,1.5403
20101229,42200,1.5403,1.5403,1.5403,1.5403
20101229,42300,1.5404,1.5404,1.5403,1.5403
20101229,42400,1.5403,1.5403,1.5403,1.5403
20101229,42500,1.5403,1.5403,1.5402,1.5402
20101229,42600,1.5403,1.5404,1.5403,1.5403
20101229,42700,1.5403,1.5403,1.5402,1.5402
20101229,42800,1.5402,1.5404,1.5401,1.5404
20101229,42900,1.5404,1.5405,1.5404,1.5404
20101229,43000,1.5405,1.5405,1.5404,1.5404
20101229,43100,1.5405,1.5405,1.5405,1.5405
20101229,43300,1.5405,1.5405,1.5404,1.5404
20101229,43400,1.5403,1.5403,1.5402,1.5403
20101229,43500,1.5403,1.5404,1.5403,1.5403
20101229,43600,1.5403,1.5403,1.5402,1.5403
20101229,43700,1.5404,1.5404,1.5403,1.5403
20101229,43800,1.5403,1.5403,1.5402,1.5403
20101229,43900,1.5403,1.5403,1.5403,1.5403
20101229,44000,1.5403,1.5403,1.5403,1.5403
20101229,44100,1.5403,1.5403,1.5403,1.5403
20101229,44200,1.5403,1.5403,1.5403,1.5403
20101229,44300,1.5403,1.5403,1.5402,1.5402
20101229,44400,1.54,1.54,1.54,1.54
20101229,44600,1.54,1.5401,1.54,1.54
20101229,44700,1.54,1.5402,1.54,1.5401
20101229,44800,1.5401,1.5401,1.5401,1.5401
20101229,44900,1.5401,1.5401,1.54,1.54
20101229,45000,1.5396,1.5396,1.5396,1.5396
20101229,45200,1.5397,1.5397,1.5397,1.5397
20101229,45400,1.5396,1.5397,1.5396,1.5397
20101229,45500,1.5397,1.5397,1.5396,1.5396
20101229,45600,1.5396,1.5396,1.5396,1.5396
20101229,45700,1.5397,1.5397,1.5397,1.5397
20101229,45800,1.5397,1.5397,1.5397,1.5397
20101229,50000,1.5397,1.5397,1.5397,1.5397
20101229,50100,1.5396,1.5396,1.5396,1.5396
20101229,50200,1.5396,1.5396,1.5395,1.5396
20101229,50300,1.5395,1.5396,1.5395,1.5395
20101229,50400,1.5395,1.5396,1.5395,1.5396
20101229,50500,1.5396,1.5396,1.5396,1.5396
20101229,50600,1.5396,1.5396,1.5396,1.5396
20101229,50700,1.5397,1.5397,1.5397,1.5397
20101229,50900,1.5397,1.5397,1.5397,1.5397
20101229,51000,1.5397,1.5397,1.5397,1.5397
20101229,51100,1.5396,1.5396,1.5396,1.5396
20101229,51300,1.5396,1.5396,1.5395,1.5396
20101229,51400,1.5397,1.5397,1.5397,1.5397
20101229,51500,1.5398,1.5398,1.5398,1.5398
20101229,51600,1.5398,1.5398,1.5398,1.5398
20101229,51800,1.5397,1.5398,1.5397,1.5397
20101229,51900,1.5396,1.5396,1.5396,1.5396
20101229,52100,1.54,1.54,1.54,1.54
20101229,52200,1.54,1.54,1.54,1.54
20101229,52400,1.5399,1.54,1.5399,1.5399
20101229,52500,1.5398,1.5398,1.5398,1.5398
20101229,52700,1.5397,1.5397,1.5397,1.5397
20101229,52800,1.5396,1.5397,1.5396,1.5397
20101229,52900,1.5397,1.5398,1.5397,1.5397
20101229,53000,1.5397,1.5397,1.5396,1.5397
20101229,53100,1.5397,1.5397,1.5397,1.5397
20101229,53200,1.5397,1.5397,1.5397,1.5397
20101229,53300,1.5397,1.5397,1.5397,1.5397
20101229,53400,1.5397,1.5397,1.5397,1.5397
20101229,53500,1.5397,1.5397,1.5396,1.5396
20101229,53600,1.5396,1.5397,1.5396,1.5397
20101229,53700,1.5396,1.5397,1.5395,1.5395
20101229,53800,1.5395,1.5396,1.5395,1.5395
20101229,53900,1.5395,1.5395,1.5395,1.5395
20101229,54000,1.5395,1.5395,1.5394,1.5394
20101229,54100,1.5388,1.5388,1.5388,1.5388
20101229,54200,1.5389,1.5389,1.5389,1.5389
20101229,54300,1.5389,1.5389,1.5389,1.5389
20101229,54500,1.5389,1.5389,1.5389,1.5389
20101229,54600,1.5391,1.5391,1.5391,1.5391
20101229,54800,1.5391,1.5391,1.5391,1.5391
20101229,54900,1.539,1.539,1.539,1.539
20101229,55000,1.539,1.539,1.539,1.539
20101229,55200,1.539,1.539,1.539,1.539
20101229,55300,1.539,1.539,1.539,1.539
20101229,55400,1.5391,1.5391,1.5391,1.5391
20101229,55600,1.5391,1.5391,1.539,1.5391
20101229,55700,1.5391,1.5391,1.5391,1.5391
20101229,55800,1.5391,1.5391,1.5391,1.5391
20101229,55900,1.539,1.539,1.539,1.539
20101229,60000,1.5382,1.5382,1.5382,1.5382
20101229,60100,1.5381,1.5381,1.5381,1.5381
20101229,60300,1.5384,1.5384,1.5384,1.5384
20101229,60500,1.5386,1.5386,1.5386,1.5386
20101229,60700,1.5384,1.5384,1.5384,1.5384
20101229,60800,1.5383,1.5383,1.5383,1.5383
20101229,60900,1.5386,1.5386,1.5386,1.5386
20101229,61000,1.5387,1.5387,1.5387,1.5387
20101229,61100,1.5386,1.5386,1.5386,1.5386
20101229,61300,1.5385,1.5386,1.5385,1.5386
20101229,61400,1.5386,1.5388,1.5386,1.5388
20101229,61500,1.5387,1.5388,1.5387,1.5387
20101229,61600,1.5386,1.5386,1.5386,1.5386
20101229,61700,1.5386,1.5386,1.5386,1.5386
20101229,61900,1.5385,1.5386,1.5385,1.5385
20101229,62000,1.5385,1.5386,1.5385,1.5386
20101229,62100,1.5386,1.5386,1.5386,1.5386
20101229,62200,1.5386,1.5386,1.5386,1.5386
20101229,62300,1.5386,1.5387,1.5386,1.5386
20101229,62400,1.5389,1.5389,1.5389,1.5389
20101229,62600,1.5388,1.5388,1.5388,1.5388
20101229,62700,1.538,1.538,1.538,1.538
20101229,62800,1.5382,1.5382,1.5382,1.5382
20101229,63000,1.5385,1.5385,1.5385,1.5385
20101229,63100,1.5385,1.5385,1.5385,1.5385
20101229,63200,1.5386,1.5386,1.5386,1.5386
20101229,63300,1.5384,1.5384,1.5384,1.5384
20101229,63500,1.5384,1.5384,1.5384,1.5384
20101229,63700,1.5384,1.5384,1.5384,1.5384
20101229,63800,1.5384,1.5384,1.5384,1.5384
20101229,63900,1.5385,1.5385,1.5385,1.5385
20101229,64000,1.5384,1.5386,1.5384,1.5386
20101229,64100,1.5386,1.5388,1.5386,1.5388
20101229,64200,1.5388,1.5389,1.5388,1.5389
20101229,64300,1.539,1.539,1.5389,1.5389
20101229,64400,1.5389,1.539,1.5389,1.5389
20101229,64500,1.5389,1.5389,1.5389,1.5389
20101229,64600,1.539,1.5394,1.539,1.5394
20101229,64700,1.5395,1.5395,1.5394,1.5394
20101229,64800,1.5395,1.5395,1.5395,1.5395
20101229,65000,1.5395,1.5395,1.5395,1.5395
20101229,65200,1.5396,1.5396,1.5396,1.5396
20101229,65400,1.5395,1.5395,1.5395,1.5395
20101229,65500,1.5395,1.5395,1.5395,1.5395
20101229,65600,1.5396,1.5396,1.5396,1.5396
20101229,65700,1.5395,1.5395,1.5395,1.5395
20101229,65800,1.5395,1.5395,1.5395,1.5395
20101229,70000,1.5396,1.5396,1.5395,1.5395
20101229,70100,1.5396,1.5396,1.5396,1.5396
20101229,70200,1.5396,1.5396,1.5396,1.5396
20101229,70300,1.5396,1.5396,1.5396,1.5396
20101229,70400,1.5395,1.5395,1.5395,1.5395
20101229,70500,1.5396,1.5396,1.5396,1.5396
20101229,70700,1.5395,1.5396,1.5395,1.5396
20101229,70800,1.5395,1.5396,1.5395,1.5395
20101229,70900,1.5395,1.5395,1.5395,1.5395
20101229,71000,1.5397,1.5397,1.5397,1.5397
20101229,71100,1.54,1.54,1.54,1.54
20101229,71200,1.5401,1.5401,1.5401,1.5401
20101229,71300,1.5402,1.5402,1.5402,1.5402
20101229,71500,1.5399,1.5399,1.5399,1.5399
20101229,71600,1.5397,1.5397,1.5397,1.5397
20101229,71800,1.5385,1.5385,1.5385,1.5385
20101229,71900,1.5387,1.5387,1.5387,1.5387
20101229,72000,1.5387,1.5387,1.5387,1.5387
20101229,72100,1.5384,1.5384,1.5384,1.5384
20101229,72200,1.5385,1.5385,1.5385,1.5385
20101229,72300,1.5386,1.5386,1.5386,1.5386
20101229,72500,1.5385,1.5386,1.5384,1.5384
20101229,72600,1.5382,1.5382,1.5382,1.5382
20101229,72700,1.5384,1.5384,1.5384,1.5384
20101229,72800,1.5385,1.5385,1.5385,1.5385
20101229,73000,1.5401,1.5401,1.5401,1.5401
20101229,73200,1.54,1.54,1.54,1.54
20101229,73300,1.5398,1.5398,1.5398,1.5398
20101229,73500,1.5399,1.5401,1.5399,1.5399
20101229,73600,1.54,1.54,1.54,1.54
20101229,73700,1.5399,1.5399,1.5399,1.5399
20101229,73900,1.5398,1.5403,1.5397,1.5403
20101229,74000,1.5401,1.5401,1.5401,1.5401
20101229,74100,1.5409,1.5409,1.5409,1.5409
20101229,74200,1.5403,1.5403,1.5403,1.5403
20101229,74400,1.5403,1.5403,1.5403,1.5403
20101229,74600,1.5402,1.5402,1.5397,1.5397
20101229,74700,1.5394,1.5394,1.5394,1.5394
20101229,74800,1.5394,1.5394,1.5394,1.5394
20101229,75000,1.5391,1.5391,1.5391,1.5391
20101229,75100,1.5388,1.5388,1.5388,1.5388
20101229,75200,1.539,1.539,1.539,1.539
20101229,75300,1.5392,1.5392,1.5392,1.5392
20101229,75400,1.5391,1.5391,1.5391,1.5391
20101229,75600,1.5397,1.5397,1.5397,1.5397
20101229,75700,1.539,1.539,1.539,1.539
20101229,75900,1.5385,1.5385,1.5385,1.5385
20101229,80000,1.538,1.538,1.538,1.538
20101229,80100,1.538,1.538,1.538,1.538
20101229,80200,1.538,1.538,1.538,1.538
20101229,80300,1.5373,1.5373,1.5373,1.5373
20101229,80400,1.5371,1.5371,1.5371,1.5371
20101229,80500,1.5361,1.5361,1.5361,1.5361
20101229,80600,1.5366,1.5366,1.5366,1.5366
20101229,80700,1.5369,1.5369,1.5369,1.5369
20101229,80900,1.537,1.5372,1.537,1.5372
20101229,81000,1.5381,1.5381,1.5381,1.5381
20101229,81100,1.5382,1.5382,1.5382,1.5382
20101229,81300,1.5381,1.5382,1.5381,1.5381
20101229,81400,1.538,1.538,1.538,1.538
20101229,81500,1.5381,1.5381,1.5381,1.5381
20101229,81600,1.5382,1.5382,1.5382,1.5382
20101229,81700,1.5382,1.5382,1.5382,1.5382
20101229,81800,1.5381,1.5381,1.5381,1.5381
20101229,81900,1.5384,1.5384,1.5384,1.5384
20101229,82100,1.5385,1.5385,1.5382,1.5382
20101229,82200,1.5384,1.5384,1.5384,1.5384
20101229,82300,1.5384,1.5384,1.5384,1.5384
20101229,82500,1.5382,1.5382,1.5382,1.5382
20101229,82600,1.5382,1.5382,1.5382,1.5382
20101229,82800,1.5382,1.5382,1.5376,1.5376
20101229,82900,1.5368,1.5368,1.5368,1.5368
20101229,83000,1.5372,1.5372,1.5372,1.5372
20101229,83100,1.5369,1.5369,1.5369,1.5369
20101229,83200,1.5371,1.5371,1.5371,1.5371
20101229,83300,1.5373,1.5373,1.5373,1.5373
20101229,83500,1.537,1.537,1.537,1.537
20101229,83600,1.5372,1.5372,1.5372,1.5372
20101229,83800,1.5369,1.5369,1.5369,1.5369
20101229,84000,1.537,1.537,1.537,1.537
20101229,84200,1.5368,1.5368,1.5368,1.5368
20101229,84300,1.5368,1.5368,1.5368,1.5368
20101229,84400,1.5369,1.5369,1.5369,1.5369
20101229,84500,1.5371,1.5371,1.5371,1.5371
20101229,84700,1.5377,1.5377,1.5377,1.5377
20101229,84800,1.5369,1.5369,1.5369,1.5369
20101229,84900,1.5369,1.5369,1.5369,1.5369
20101229,85100,1.5372,1.5372,1.5372,1.5372
20101229,85200,1.5372,1.5372,1.5372,1.5372
20101229,85400,1.5372,1.5372,1.5372,1.5372
20101229,85500,1.5372,1.5372,1.5372,1.5372
20101229,85700,1.5379,1.5379,1.5379,1.5379
20101229,85900,1.538,1.538,1.538,1.538
20101229,90000,1.5381,1.5381,1.5381,1.5381
20101229,90200,1.5382,1.5382,1.5382,1.5382
20101229,90300,1.538,1.538,1.538,1.538
20101229,90400,1.5379,1.5379,1.5379,1.5379
20101229,90500,1.5371,1.5371,1.5371,1.5371
20101229,90700,1.5371,1.5372,1.5369,1.5369
20101229,90800,1.5369,1.5369,1.5367,1.5368
20101229,90900,1.5369,1.5375,1.5369,1.5375
20101229,91000,1.5376,1.5376,1.5371,1.5373
20101229,91100,1.5383,1.5383,1.5383,1.5383
20101229,91200,1.5383,1.5383,1.5383,1.5383
20101229,91400,1.5383,1.5383,1.5382,1.5383
20101229,91500,1.5383,1.5383,1.5383,1.5383
20101229,91700,1.5384,1.5385,1.5382,1.5382
20101229,91800,1.5381,1.5383,1.5381,1.5383
20101229,91900,1.5382,1.5382,1.5382,1.5382
20101229,92100,1.5388,1.5388,1.5388,1.5388
20101229,92200,1.5387,1.5387,1.5387,1.5387
20101229,92300,1.5386,1.5386,1.5386,1.5386
20101229,92400,1.5386,1.5386,1.5386,1.5386
20101229,92600,1.5386,1.5386,1.5386,1.5386
20101229,92800,1.5387,1.5387,1.5387,1.5387
20101229,92900,1.5385,1.5385,1.5385,1.5385
20101229,93000,1.5385,1.5385,1.5385,1.5385
20101229,93200,1.5383,1.5383,1.5383,1.5383
20101229,93300,1.538,1.538,1.538,1.538
20101229,93400,1.538,1.538,1.538,1.538
20101229,93600,1.5381,1.5381,1.5378,1.5378
20101229,93700,1.5379,1.5383,1.5379,1.5383
20101229,93800,1.5382,1.5382,1.5381,1.5381
20101229,93900,1.5382,1.5385,1.538,1.5384
20101229,94000,1.5385,1.5385,1.5383,1.5383
20101229,94100,1.5381,1.5381,1.5381,1.5381
20101229,94200,1.5381,1.5381,1.5381,1.5381
20101229,94400,1.5384,1.5384,1.5384,1.5384
20101229,94600,1.5383,1.5383,1.5382,1.5382
20101229,94700,1.5383,1.5387,1.5383,1.5385
20101229,94800,1.5384,1.5386,1.5382,1.5383
20101229,94900,1.5383,1.5383,1.5383,1.5383
20101229,95000,1.5383,1.5383,1.5383,1.5383
20101229,95100,1.5379,1.5379,1.5379,1.5379
20101229,95200,1.5378,1.5378,1.5378,1.5378
20101229,95400,1.5376,1.5376,1.5376,1.5376
20101229,95600,1.5377,1.5377,1.5375,1.5376
20101229,95700,1.5375,1.5376,1.5374,1.5374
20101229,95800,1.5374,1.5375,1.5374,1.5375
20101229,95900,1.5369,1.5369,1.5369,1.5369
20101229,100000,1.5374,1.5374,1.5374,1.5374
20101229,100200,1.5373,1.5373,1.5372,1.5372
20101229,100300,1.5373,1.5373,1.5368,1.5369
20101229,100400,1.537,1.5371,1.537,1.5371
20101229,100500,1.537,1.537,1.5367,1.537
20101229,100600,1.537,1.5372,1.537,1.5371
20101229,100700,1.5374,1.5374,1.5374,1.5374
20101229,100800,1.5377,1.5377,1.5377,1.5377
20101229,101000,1.5381,1.5381,1.5381,1.5381
20101229,101100,1.5382,1.5382,1.5382,1.5382
20101229,101300,1.5381,1.5381,1.5379,1.5379
20101229,101400,1.5381,1.5381,1.5381,1.5381
20101229,101500,1.5382,1.5382,1.5382,1.5382
20101229,101700,1.5383,1.5385,1.5382,1.5384
20101229,101800,1.5385,1.5385,1.5384,1.5384
20101229,101900,1.5384,1.5384,1.5384,1.5384
20101229,102100,1.5381,1.5381,1.5381,1.5381
20101229,102300,1.538,1.538,1.538,1.538
20101229,102500,1.5379,1.5379,1.5378,1.5378
20101229,102600,1.5377,1.5379,1.5377,1.5379
20101229,102700,1.5379,1.538,1.5379,1.538
20101229,102800,1.5376,1.5376,1.5376,1.5376
20101229,102900,1.5375,1.5375,1.5375,1.5375
20101229,103000,1.5373,1.5373,1.5373,1.5373
20101229,103100,1.5371,1.5371,1.5371,1.5371
20101229,103200,1.5374,1.5374,1.5374,1.5374
20101229,103300,1.5373,1.5373,1.5373,1.5373
20101229,103500,1.5379,1.5379,1.5379,1.5379
20101229,103600,1.5377,1.5377,1.5377,1.5377
20101229,103800,1.5378,1.5379,1.5375,1.5379
20101229,103900,1.5378,1.5378,1.5376,1.5376
20101229,104000,1.5376,1.5376,1.5375,1.5375
20101229,104100,1.5376,1.5376,1.5372,1.5376
20101229,104200,1.5372,1.5372,1.5372,1.5372
20101229,104400,1.5377,1.5377,1.5377,1.5377
20101229,104600,1.5379,1.5379,1.5379,1.5379
20101229,104800,1.5378,1.5378,1.5376,1.5376
20101229,104900,1.5375,1.5379,1.5375,1.5376
20101229,105000,1.5376,1.5376,1.5375,1.5376
20101229,105100,1.5375,1.5381,1.5375,1.5381
20101229,105200,1.538,1.5385,1.538,1.5384
20101229,105300,1.5384,1.5384,1.5384,1.5384
20101229,105400,1.5391,1.5391,1.5391,1.5391
20101229,105500,1.539,1.539,1.539,1.539
20101229,105600,1.5395,1.5395,1.5395,1.5395
20101229,105700,1.5387,1.5387,1.5387,1.5387
20101229,105800,1.539,1.539,1.539,1.539
20101229,105900,1.5397,1.5397,1.5397,1.5397
20101229,110000,1.5397,1.5397,1.5397,1.5397
20101229,110100,1.5395,1.5395,1.5395,1.5395
20101229,110300,1.5391,1.5391,1.5391,1.5391
20101229,110500,1.5394,1.5394,1.5394,1.5394
20101229,110600,1.5392,1.5392,1.5392,1.5392
20101229,110800,1.539,1.539,1.539,1.539
20101229,110900,1.5387,1.5387,1.5387,1.5387
20101229,111100,1.5388,1.5388,1.5388,1.5388
20101229,111200,1.5389,1.5389,1.5389,1.5389
20101229,111400,1.5388,1.5388,1.5388,1.5388
20101229,111600,1.5387,1.5389,1.5386,1.5386
20101229,111700,1.5385,1.5385,1.5385,1.5385
20101229,111800,1.5384,1.5384,1.5384,1.5384
20101229,112000,1.5382,1.5382,1.5382,1.5382
20101229,112100,1.5383,1.5383,1.5383,1.5383
20101229,112200,1.538,1.538,1.538,1.538
20101229,112400,1.5384,1.5384,1.5384,1.5384
20101229,112600,1.5382,1.5382,1.5382,1.5382
20101229,112700,1.5381,1.5381,1.5381,1.5381
20101229,112900,1.5384,1.5384,1.5384,1.5384
20101229,113000,1.5391,1.5391,1.5391,1.5391
20101229,113100,1.539,1.539,1.539,1.539
20101229,113200,1.5391,1.5391,1.5391,1.5391
20101229,113300,1.5393,1.5393,1.5393,1.5393
20101229,113400,1.5389,1.5389,1.5389,1.5389
20101229,113500,1.539,1.539,1.539,1.539
20101229,113700,1.5382,1.5382,1.5382,1.5382
20101229,113800,1.5384,1.5384,1.5384,1.5384
20101229,114000,1.5384,1.5385,1.5383,1.5384
20101229,114100,1.5386,1.5386,1.5386,1.5386
20101229,114200,1.5386,1.5386,1.5386,1.5386
20101229,114300,1.5386,1.5386,1.5386,1.5386
20101229,114400,1.5386,1.5386,1.5386,1.5386
20101229,114500,1.5391,1.5391,1.5391,1.5391
20101229,114600,1.5391,1.5391,1.5391,1.5391
20101229,114700,1.5393,1.5393,1.5393,1.5393
20101229,114900,1.5391,1.5391,1.5391,1.5391
20101229,115000,1.5389,1.5389,1.5389,1.5389
20101229,115200,1.5396,1.5396,1.5396,1.5396
20101229,115400,1.5394,1.5394,1.5394,1.5394
20101229,115600,1.5392,1.5392,1.5392,1.5392
20101229,115800,1.5392,1.5392,1.5392,1.5392
20101229,120000,1.5393,1.5393,1.5393,1.5393
20101229,120100,1.5396,1.5396,1.5396,1.5396
20101229,120300,1.5401,1.5401,1.5401,1.5401
20101229,120400,1.54,1.54,1.54,1.54
20101229,120500,1.54,1.54,1.54,1.54
20101229,120600,1.5393,1.5393,1.5393,1.5393
20101229,120700,1.5391,1.5391,1.5391,1.5391
20101229,120800,1.5394,1.5394,1.5394,1.5394
20101229,120900,1.5396,1.5396,1.5396,1.5396
20101229,121100,1.5393,1.5393,1.5393,1.5393
20101229,121200,1.5396,1.5396,1.5396,1.5396
20101229,121300,1.5395,1.5395,1.5395,1.5395
20101229,121500,1.5388,1.5388,1.5388,1.5388
20101229,121600,1.5389,1.5389,1.5389,1.5389
20101229,121700,1.5384,1.5384,1.5384,1.5384
20101229,121800,1.5381,1.5381,1.5381,1.5381
20101229,121900,1.5386,1.5386,1.5386,1.5386
20101229,122000,1.5391,1.5391,1.5391,1.5391
20101229,122100,1.5386,1.5386,1.5386,1.5386
20101229,122200,1.5386,1.5386,1.5386,1.5386
20101229,122300,1.5387,1.5387,1.5387,1.5387
20101229,122500,1.5387,1.5387,1.5387,1.5387
20101229,122600,1.5386,1.5386,1.5386,1.5386
20101229,122800,1.5392,1.5392,1.5392,1.5392
20101229,122900,1.5398,1.5398,1.5398,1.5398
20101229,123000,1.5393,1.5393,1.5393,1.5393
20101229,123100,1.5394,1.5394,1.5394,1.5394
20101229,123200,1.5393,1.5393,1.5393,1.5393
20101229,123300,1.5394,1.5394,1.5394,1.5394
20101229,123400,1.5395,1.5395,1.5395,1.5395
20101229,123600,1.5392,1.5392,1.5392,1.5392
20101229,123700,1.539,1.539,1.539,1.539
20101229,123900,1.539,1.5392,1.539,1.5391
20101229,124000,1.5396,1.5396,1.5396,1.5396
20101229,124100,1.5397,1.5397,1.5397,1.5397
20101229,124200,1.5394,1.5394,1.5394,1.5394
20101229,124300,1.5392,1.5392,1.5392,1.5392
20101229,124400,1.5389,1.5389,1.5389,1.5389
20101229,124600,1.539,1.539,1.539,1.539
20101229,124800,1.5388,1.5388,1.5388,1.5388
20101229,124900,1.5387,1.5387,1.5387,1.5387
20101229,125000,1.5389,1.5389,1.5389,1.5389
20101229,125100,1.539,1.539,1.539,1.539
20101229,125300,1.5387,1.5387,1.5387,1.5387
20101229,125400,1.5389,1.5389,1.5389,1.5389
20101229,125500,1.539,1.539,1.539,1.539
20101229,125600,1.539,1.539,1.539,1.539
20101229,125800,1.5381,1.5381,1.5381,1.5381
20101229,125900,1.5373,1.5373,1.5373,1.5373
20101229,130000,1.5377,1.5377,1.5377,1.5377
20101229,130100,1.5375,1.5375,1.5375,1.5375
20101229,130300,1.5372,1.5372,1.5372,1.5372
20101229,130400,1.5374,1.5374,1.5374,1.5374
20101229,130600,1.5375,1.5375,1.5375,1.5375
20101229,130700,1.5378,1.5378,1.5378,1.5378
20101229,130900,1.5378,1.538,1.5378,1.538
20101229,131000,1.5379,1.538,1.5377,1.538
20101229,131100,1.5379,1.5379,1.5379,1.5379
20101229,131200,1.5379,1.5379,1.5379,1.5379
20101229,131400,1.5376,1.5376,1.5376,1.5376
20101229,131500,1.5381,1.5381,1.5381,1.5381
20101229,131600,1.5379,1.5379,1.5379,1.5379
20101229,131700,1.5379,1.5379,1.5379,1.5379
20101229,131800,1.5379,1.5379,1.5379,1.5379
20101229,131900,1.5376,1.5376,1.5376,1.5376
20101229,132000,1.5373,1.5373,1.5373,1.5373
20101229,132100,1.5376,1.5376,1.5376,1.5376
20101229,132300,1.5375,1.5375,1.5372,1.5374
20101229,132400,1.5373,1.5374,1.5373,1.5374
20101229,132500,1.5371,1.5371,1.5371,1.5371
20101229,132700,1.5375,1.5375,1.5375,1.5375
20101229,132900,1.5381,1.5381,1.5381,1.5381
20101229,133100,1.5384,1.5384,1.5384,1.5384
20101229,133200,1.5383,1.5383,1.5383,1.5383
20101229,133300,1.5386,1.5386,1.5386,1.5386
20101229,133500,1.539,1.539,1.539,1.539
20101229,133600,1.5389,1.5389,1.5389,1.5389
20101229,133700,1.5385,1.5385,1.5385,1.5385
20101229,133800,1.5387,1.5387,1.5387,1.5387
20101229,133900,1.5386,1.5386,1.5386,1.5386
20101229,134000,1.5388,1.5388,1.5388,1.5388
20101229,134200,1.5389,1.5389,1.5385,1.5385
20101229,134300,1.5384,1.5384,1.5384,1.5384
20101229,134500,1.5384,1.5385,1.5384,1.5385
20101229,134600,1.5387,1.5387,1.5387,1.5387
20101229,134800,1.5388,1.5388,1.5388,1.5388
20101229,134900,1.5387,1.5387,1.5387,1.5387
20101229,135000,1.5385,1.5385,1.5385,1.5385
20101229,135200,1.5386,1.5386,1.5383,1.5385
20101229,135300,1.5388,1.5388,1.5388,1.5388
20101229,135500,1.539,1.539,1.539,1.539
20101229,135600,1.5388,1.5388,1.5388,1.5388
20101229,135700,1.539,1.539,1.539,1.539
20101229,135800,1.5391,1.5391,1.5391,1.5391
20101229,135900,1.5393,1.5393,1.5393,1.5393
20101229,140000,1.5397,1.5397,1.5397,1.5397
20101229,140100,1.5396,1.5396,1.5396,1.5396
20101229,140300,1.5391,1.5391,1.5391,1.5391
20101229,140500,1.539,1.539,1.539,1.539
20101229,140600,1.539,1.539,1.539,1.539
20101229,140700,1.5395,1.5395,1.5395,1.5395
20101229,140900,1.5396,1.5397,1.5394,1.5397
20101229,141000,1.5398,1.5398,1.5395,1.5395
20101229,141100,1.5396,1.5396,1.5396,1.5396
20101229,141200,1.5397,1.5397,1.5397,1.5397
20101229,141300,1.5395,1.5395,1.5395,1.5395
20101229,141500,1.5396,1.5396,1.5396,1.5396
20101229,141600,1.5397,1.5397,1.5397,1.5397
20101229,141700,1.5398,1.5398,1.5398,1.5398
20101229,141800,1.5398,1.5398,1.5398,1.5398
20101229,141900,1.5398,1.5398,1.5398,1.5398
20101229,142100,1.5402,1.5402,1.5402,1.5402
20101229,142200,1.54,1.54,1.54,1.54
20101229,142400,1.5402,1.5402,1.5402,1.5402
20101229,142500,1.5408,1.5408,1.5408,1.5408
20101229,142600,1.5409,1.5409,1.5409,1.5409
20101229,142700,1.5416,1.5416,1.5416,1.5416
20101229,142800,1.5415,1.5415,1.5415,1.5415
20101229,142900,1.5415,1.5415,1.5415,1.5415
20101229,143100,1.5416,1.5416,1.5416,1.5416
20101229,143200,1.542,1.542,1.542,1.542
20101229,143400,1.5421,1.5422,1.5421,1.5422
20101229,143500,1.5432,1.5432,1.5432,1.5432
20101229,143600,1.5441,1.5441,1.5441,1.5441
20101229,143700,1.5437,1.5437,1.5437,1.5437
20101229,143900,1.5436,1.5436,1.5436,1.5436
20101229,144100,1.5444,1.5444,1.5444,1.5444
20101229,144200,1.5443,1.5443,1.5443,1.5443
20101229,144400,1.5437,1.5437,1.5437,1.5437
20101229,144500,1.5439,1.5439,1.5439,1.5439
20101229,144600,1.5439,1.5439,1.5439,1.5439
20101229,144700,1.5439,1.5439,1.5439,1.5439
20101229,144800,1.5441,1.5441,1.5441,1.5441
20101229,144900,1.5439,1.5439,1.5439,1.5439
20101229,145000,1.5438,1.5438,1.5438,1.5438
20101229,145100,1.5434,1.5434,1.5434,1.5434
20101229,145200,1.5437,1.5437,1.5437,1.5437
20101229,145400,1.5436,1.5436,1.5436,1.5436
20101229,145500,1.5432,1.5432,1.5432,1.5432
20101229,145700,1.5433,1.5433,1.5431,1.5432
20101229,145800,1.5428,1.5428,1.5428,1.5428
20101229,145900,1.5429,1.5429,1.5429,1.5429
20101229,150000,1.5432,1.5432,1.5432,1.5432
20101229,150200,1.5433,1.5433,1.5433,1.5433
20101229,150300,1.5433,1.5433,1.5433,1.5433
20101229,150400,1.5433,1.5433,1.5433,1.5433
20101229,150500,1.5433,1.5433,1.5433,1.5433
20101229,150600,1.5429,1.5429,1.5429,1.5429
20101229,150700,1.5432,1.5432,1.5432,1.5432
20101229,150900,1.5427,1.5427,1.5427,1.5427
20101229,151000,1.5427,1.5427,1.5427,1.5427
20101229,151200,1.5428,1.5429,1.5428,1.5428
20101229,151300,1.5431,1.5431,1.5431,1.5431
20101229,151400,1.5437,1.5437,1.5437,1.5437
20101229,151600,1.5438,1.5438,1.5438,1.5438
20101229,151800,1.5437,1.5438,1.5432,1.5437
20101229,151900,1.5443,1.5443,1.5443,1.5443
20101229,152000,1.544,1.544,1.544,1.544
20101229,152200,1.5441,1.5441,1.5439,1.5439
20101229,152300,1.5437,1.5437,1.5437,1.5437
20101229,152500,1.544,1.544,1.544,1.544
20101229,152600,1.5437,1.5437,1.5437,1.5437
20101229,152800,1.5436,1.5436,1.5436,1.5436
20101229,152900,1.5438,1.5438,1.5438,1.5438
20101229,153000,1.5436,1.5436,1.5436,1.5436
20101229,153200,1.5433,1.5433,1.5433,1.5433
20101229,153300,1.5433,1.5433,1.5433,1.5433
20101229,153500,1.5433,1.5433,1.5433,1.5433
20101229,153600,1.5431,1.5431,1.5431,1.5431
20101229,153700,1.5429,1.5429,1.5429,1.5429
20101229,153800,1.5428,1.5428,1.5428,1.5428
20101229,153900,1.5426,1.5426,1.5426,1.5426
20101229,154100,1.5427,1.543,1.5426,1.543
20101229,154200,1.5429,1.5429,1.5429,1.5429
20101229,154300,1.543,1.543,1.543,1.543
20101229,154500,1.5433,1.5433,1.5433,1.5433
20101229,154700,1.5432,1.5432,1.5432,1.5432
20101229,154800,1.5432,1.5432,1.5432,1.5432
20101229,154900,1.5432,1.5432,1.5432,1.5432
20101229,155000,1.5437,1.5437,1.5437,1.5437
20101229,155200,1.5438,1.5438,1.5438,1.5438
20101229,155300,1.5437,1.5437,1.5437,1.5437
20101229,155500,1.5438,1.5438,1.5437,1.5437
20101229,155600,1.5435,1.5435,1.5435,1.5435
20101229,155800,1.5434,1.5434,1.5434,1.5434
20101229,155900,1.5421,1.5421,1.5421,1.5421
20101229,160000,1.5424,1.5424,1.5424,1.5424
20101229,160200,1.5429,1.5429,1.5429,1.5429
20101229,160300,1.5432,1.5432,1.5432,1.5432
20101229,160500,1.5432,1.5433,1.5432,1.5432
20101229,160600,1.5431,1.5431,1.5431,1.5431
20101229,160700,1.543,1.543,1.543,1.543
20101229,160900,1.5431,1.5432,1.543,1.5431
20101229,161000,1.5431,1.5431,1.5429,1.543
20101229,161100,1.5429,1.5429,1.5429,1.5429
20101229,161300,1.543,1.5432,1.5429,1.543
20101229,161400,1.5428,1.5428,1.5428,1.5428
20101229,161500,1.5432,1.5432,1.5432,1.5432
20101229,161600,1.5433,1.5433,1.5433,1.5433
20101229,161800,1.5433,1.5433,1.5431,1.5432
20101229,161900,1.5431,1.5431,1.5431,1.5431
20101229,162000,1.5431,1.5431,1.5431,1.5431
20101229,162100,1.5431,1.5431,1.5431,1.5431
20101229,162200,1.5434,1.5434,1.5434,1.5434
20101229,162300,1.5435,1.5435,1.5435,1.5435
20101229,162400,1.5434,1.5434,1.5434,1.5434
20101229,162500,1.5435,1.5435,1.5435,1.5435
20101229,162700,1.5436,1.5436,1.5436,1.5436
20101229,162800,1.5436,1.5436,1.5436,1.5436
20101229,163000,1.5436,1.5436,1.5435,1.5435
20101229,163100,1.5435,1.5435,1.5435,1.5435
20101229,163300,1.5434,1.5434,1.5434,1.5434
20101229,163400,1.5439,1.5439,1.5439,1.5439
20101229,163500,1.544,1.5442,1.544,1.544
20101229,163600,1.5443,1.5443,1.5443,1.5443
20101229,163700,1.5443,1.5443,1.5443,1.5443
20101229,163800,1.5448,1.5448,1.5448,1.5448
20101229,163900,1.5448,1.5448,1.5448,1.5448
20101229,164000,1.5448,1.5448,1.5448,1.5448
20101229,164100,1.5448,1.5448,1.5448,1.5448
20101229,164300,1.5447,1.5447,1.5447,1.5447
20101229,164400,1.5442,1.5442,1.5442,1.5442
20101229,164500,1.5452,1.5452,1.5452,1.5452
20101229,164600,1.5452,1.5452,1.5452,1.5452
20101229,164700,1.5453,1.5453,1.5453,1.5453
20101229,164900,1.5454,1.5455,1.5453,1.5455
20101229,165000,1.5457,1.5457,1.5457,1.5457
20101229,165100,1.5456,1.5456,1.5456,1.5456
20101229,165200,1.5459,1.5459,1.5459,1.5459
20101229,165300,1.546,1.546,1.546,1.546
20101229,165500,1.5457,1.5457,1.5457,1.5457
20101229,165600,1.5456,1.5456,1.5456,1.5456
20101229,165800,1.5456,1.5456,1.5456,1.5456
20101229,165900,1.5458,1.5458,1.5458,1.5458
20101229,170000,1.546,1.546,1.546,1.546
20101229,170100,1.5462,1.5462,1.5462,1.5462
20101229,170200,1.5463,1.5463,1.5462,1.5463
20101229,170400,1.5462,1.5462,1.5461,1.5461
20101229,170500,1.5464,1.5464,1.5464,1.5464
20101229,170700,1.5463,1.5464,1.5462,1.5462
20101229,170800,1.5463,1.5463,1.5463,1.5463
20101229,170900,1.5461,1.5461,1.5461,1.5461
20101229,171000,1.5457,1.5457,1.5457,1.5457
20101229,171100,1.5458,1.5458,1.5458,1.5458
20101229,171200,1.5458,1.5458,1.5458,1.5458
20101229,171400,1.5458,1.5458,1.5457,1.5457
20101229,171500,1.5457,1.5457,1.5455,1.5456
20101229,171600,1.5458,1.5458,1.5458,1.5458
20101229,171700,1.546,1.546,1.546,1.546
20101229,171800,1.5461,1.5461,1.5461,1.5461
20101229,172000,1.546,1.546,1.546,1.546
20101229,172200,1.5461,1.5461,1.5459,1.546
20101229,172300,1.5462,1.5462,1.5462,1.5462
20101229,172400,1.5463,1.5463,1.5463,1.5463
20101229,172600,1.5462,1.5462,1.5462,1.5462
20101229,172700,1.5462,1.5462,1.5462,1.5462
20101229,172800,1.5461,1.5461,1.5461,1.5461
20101229,172900,1.546,1.546,1.5458,1.546
20101229,173100,1.5458,1.5458,1.5458,1.5458
20101229,173200,1.546,1.546,1.546,1.546
20101229,173400,1.5461,1.5461,1.5461,1.5461
20101229,173500,1.5461,1.5461,1.5461,1.5461
20101229,173600,1.546,1.546,1.546,1.546
20101229,173700,1.546,1.546,1.546,1.546
20101229,173900,1.546,1.546,1.5459,1.5459
20101229,174000,1.5458,1.5458,1.5458,1.5458
20101229,174100,1.5458,1.5458,1.5458,1.5458
20101229,174200,1.5457,1.5457,1.5457,1.5457
20101229,174400,1.5459,1.5459,1.5459,1.5459
20101229,174500,1.5458,1.546,1.5458,1.5459
20101229,174600,1.5462,1.5462,1.5462,1.5462
20101229,174800,1.5462,1.5465,1.5461,1.5461
20101229,174900,1.5461,1.5463,1.5461,1.5463
20101229,175000,1.5463,1.5463,1.5462,1.5462
20101229,175100,1.5463,1.5463,1.5463,1.5463
20101229,175300,1.5464,1.5464,1.5464,1.5464
20101229,175400,1.5466,1.5466,1.5466,1.5466
20101229,175600,1.5466,1.5467,1.5465,1.5467
20101229,175700,1.548,1.548,1.548,1.548
20101229,175900,1.5482,1.5482,1.5482,1.5482
20101229,180000,1.5488,1.5489,1.5482,1.5482
20101229,180100,1.5481,1.5483,1.548,1.548
20101229,180200,1.5481,1.5486,1.5481,1.5485
20101229,180300,1.5486,1.5494,1.5486,1.5491
20101229,180400,1.5491,1.5497,1.5491,1.5497
20101229,180500,1.5496,1.5496,1.5492,1.5493
20101229,180600,1.5494,1.5503,1.5494,1.55
20101229,180700,1.5499,1.5499,1.5496,1.5496
20101229,180800,1.5495,1.5495,1.5493,1.5494
20101229,180900,1.5493,1.5496,1.5493,1.5496
20101229,181000,1.5495,1.5495,1.5492,1.5494
20101229,181100,1.5493,1.5493,1.549,1.5492
20101229,181200,1.5493,1.5493,1.549,1.5491
20101229,181300,1.549,1.5491,1.549,1.549
20101229,181400,1.549,1.549,1.5489,1.549
20101229,181500,1.549,1.549,1.5489,1.549
20101229,181600,1.5491,1.5494,1.5491,1.5494
20101229,181700,1.5495,1.5499,1.5495,1.5498
20101229,181800,1.5498,1.5498,1.5496,1.5497
20101229,181900,1.5497,1.55,1.5496,1.5499
20101229,182000,1.5498,1.5498,1.5497,1.5497
20101229,182100,1.5497,1.5499,1.5497,1.5498
20101229,182200,1.5499,1.55,1.5498,1.55
20101229,182300,1.5501,1.5504,1.55,1.5504
20101229,182400,1.5505,1.5505,1.5503,1.5504
20101229,182500,1.5504,1.5508,1.5504,1.5508
20101229,182600,1.5507,1.5508,1.5501,1.5501
20101229,182700,1.55,1.5501,1.55,1.55
20101229,182800,1.55,1.55,1.5499,1.55
20101229,182900,1.55,1.55,1.5499,1.55
20101229,183000,1.5499,1.5499,1.5497,1.5497
20101229,183100,1.5498,1.5498,1.5498,1.5498
20101229,183200,1.5498,1.5499,1.5498,1.5498
20101229,183300,1.5497,1.5498,1.5497,1.5497
20101229,183400,1.5497,1.5498,1.5496,1.5497
20101229,183500,1.5497,1.5497,1.5495,1.5495
20101229,183600,1.5494,1.5494,1.5493,1.5493
20101229,183700,1.5494,1.5494,1.5493,1.5494
20101229,183800,1.5493,1.5493,1.5492,1.5493
20101229,183900,1.5494,1.5494,1.5493,1.5494
20101229,184000,1.5493,1.5493,1.5489,1.5489
20101229,184100,1.5488,1.5489,1.5488,1.5489
20101229,184200,1.5489,1.549,1.5489,1.549
20101229,184300,1.549,1.549,1.5489,1.549
20101229,184400,1.5491,1.5498,1.5491,1.5495
20101229,184500,1.5494,1.5495,1.5494,1.5495
20101229,184600,1.5496,1.5496,1.5495,1.5495
20101229,184700,1.5496,1.5498,1.5495,1.5497
20101229,184800,1.5496,1.5496,1.5496,1.5496
20101229,184900,1.5497,1.5499,1.5497,1.5498
20101229,185000,1.5497,1.5497,1.5494,1.5495
20101229,185100,1.5495,1.5495,1.5495,1.5495
20101229,185200,1.5495,1.5498,1.5495,1.5497
20101229,185300,1.5497,1.5499,1.5497,1.5499
20101229,185400,1.55,1.55,1.5497,1.5498
20101229,185500,1.5499,1.5499,1.5497,1.5497
20101229,185600,1.5497,1.5497,1.5495,1.5496
20101229,185700,1.5496,1.5496,1.5495,1.5496
20101229,185800,1.5495,1.5496,1.5495,1.5495
20101229,185900,1.5495,1.5495,1.5492,1.5492
20101229,190000,1.5493,1.5493,1.5493,1.5493
20101229,190100,1.5494,1.5494,1.5493,1.5494
20101229,190200,1.5494,1.5494,1.5494,1.5494
20101229,190300,1.5494,1.5494,1.5494,1.5494
20101229,190400,1.5494,1.5494,1.5494,1.5494
20101229,190500,1.5493,1.5493,1.5493,1.5493
20101229,190600,1.5493,1.5494,1.5493,1.5493
20101229,190700,1.5493,1.5494,1.5493,1.5494
20101229,190800,1.5494,1.5495,1.5494,1.5495
20101229,190900,1.5494,1.5498,1.5494,1.5498
20101229,191000,1.55,1.55,1.5497,1.5497
20101229,191100,1.5498,1.5498,1.5497,1.5498
20101229,191200,1.5498,1.5499,1.5497,1.5498
20101229,191300,1.5499,1.5501,1.5499,1.5501
20101229,191400,1.55,1.5501,1.55,1.55
20101229,191500,1.55,1.55,1.5497,1.5497
20101229,191600,1.5498,1.5502,1.5498,1.55
20101229,191700,1.5501,1.5501,1.55,1.5501
20101229,191800,1.5501,1.5501,1.55,1.55
20101229,191900,1.5501,1.5501,1.5498,1.5499
20101229,192000,1.5499,1.5499,1.5498,1.5498
20101229,192100,1.5497,1.5499,1.5497,1.5498
20101229,192200,1.5497,1.5498,1.5497,1.5498
20101229,192300,1.5498,1.5498,1.5495,1.5495
20101229,192400,1.5496,1.5496,1.5496,1.5496
20101229,192500,1.5496,1.5496,1.5496,1.5496
20101229,192600,1.5496,1.5496,1.5496,1.5496
20101229,192700,1.5496,1.55,1.5496,1.55
20101229,192800,1.5499,1.5499,1.5495,1.5495
20101229,192900,1.5496,1.5496,1.5495,1.5496
20101229,193000,1.5496,1.5497,1.5496,1.5497
20101229,193100,1.5497,1.5498,1.5497,1.5498
20101229,193200,1.5498,1.5499,1.5498,1.5499
20101229,193300,1.5498,1.55,1.5498,1.5499
20101229,193400,1.55,1.5502,1.55,1.55
20101229,193500,1.55,1.55,1.5499,1.55
20101229,193600,1.55,1.55,1.55,1.55
20101229,193700,1.5499,1.5499,1.5498,1.5499
20101229,193800,1.5499,1.5499,1.5498,1.5498
20101229,193900,1.5498,1.5499,1.5498,1.5499
20101229,194000,1.55,1.5501,1.5497,1.5497
20101229,194100,1.5497,1.5498,1.5497,1.5498
20101229,194200,1.5498,1.5498,1.5497,1.5497
20101229,194300,1.5497,1.5497,1.5496,1.5497
20101229,194400,1.5497,1.5497,1.5495,1.5497
20101229,194500,1.5497,1.5498,1.5496,1.5498
20101229,194600,1.5498,1.5498,1.5496,1.5497
20101229,194700,1.5497,1.5497,1.5497,1.5497
20101229,194800,1.5497,1.5502,1.5497,1.5501
20101229,194900,1.55,1.5501,1.55,1.55
20101229,195000,1.5499,1.5499,1.5498,1.5499
20101229,195100,1.5498,1.5498,1.5498,1.5498
20101229,195200,1.5498,1.5499,1.5498,1.5499
20101229,195300,1.5499,1.5499,1.5498,1.5498
20101229,195400,1.5498,1.55,1.5498,1.5499
20101229,195500,1.55,1.55,1.5499,1.5499
20101229,195600,1.5499,1.5502,1.5499,1.5502
20101229,195700,1.5501,1.5502,1.5501,1.5502
20101229,195800,1.5501,1.5502,1.5501,1.5502
20101229,195900,1.5503,1.5505,1.5503,1.5505
20101229,200000,1.5504,1.5508,1.5504,1.5507
20101229,200100,1.5505,1.5508,1.5505,1.5505
20101229,200200,1.5505,1.5507,1.5505,1.5506
20101229,200300,1.5506,1.5506,1.5501,1.5501
20101229,200400,1.5502,1.5503,1.5501,1.5503
20101229,200500,1.5503,1.5503,1.5502,1.5503
20101229,200600,1.5503,1.5504,1.5503,1.5503
20101229,200700,1.5504,1.5505,1.5504,1.5505
20101229,200800,1.5506,1.5507,1.5506,1.5506
20101229,200900,1.5505,1.5509,1.5505,1.5509
20101229,201000,1.551,1.5512,1.5509,1.5512
20101229,201100,1.5512,1.5513,1.5512,1.5513
20101229,201200,1.5513,1.5515,1.5513,1.5515
20101229,201300,1.5515,1.5515,1.5513,1.5513
20101229,201400,1.5513,1.5514,1.5513,1.5513
20101229,201500,1.5513,1.5514,1.5513,1.5514
20101229,201600,1.5514,1.5514,1.5513,1.5514
20101229,201700,1.5515,1.5516,1.5515,1.5515
20101229,201800,1.5514,1.5514,1.5512,1.5513
20101229,201900,1.5513,1.5514,1.5513,1.5514
20101229,202000,1.5513,1.5513,1.5512,1.5512
20101229,202100,1.5512,1.5513,1.5512,1.5512
20101229,202200,1.5513,1.5513,1.5512,1.5512
20101229,202300,1.5512,1.5512,1.5511,1.5511
20101229,202400,1.5511,1.5512,1.551,1.5511
20101229,202500,1.5511,1.5511,1.551,1.551
20101229,202600,1.551,1.551,1.5508,1.5508
20101229,202700,1.5508,1.5508,1.5508,1.5508
20101229,202800,1.5508,1.5508,1.5508,1.5508
20101229,202900,1.5508,1.551,1.5508,1.5508
20101229,203000,1.5508,1.5508,1.5508,1.5508
20101229,203100,1.5508,1.5508,1.5507,1.5508
20101229,203200,1.5509,1.5511,1.5507,1.5507
20101229,203300,1.5506,1.5506,1.55,1.55
20101229,203400,1.5501,1.5504,1.5501,1.5502
20101229,203500,1.5501,1.5503,1.5501,1.5503
20101229,203600,1.5503,1.5504,1.5503,1.5503
20101229,203700,1.5502,1.5503,1.5502,1.5503
20101229,203800,1.5504,1.5506,1.5503,1.5506
20101229,203900,1.5505,1.5508,1.5505,1.5507
20101229,204000,1.5508,1.5509,1.5506,1.5507
20101229,204100,1.5508,1.5508,1.5505,1.5505
20101229,204200,1.5504,1.5504,1.5501,1.5501
20101229,204300,1.5502,1.5502,1.5502,1.5502
20101229,204400,1.5502,1.5503,1.5501,1.5503
20101229,204500,1.5503,1.5503,1.5503,1.5503
20101229,204600,1.5504,1.5504,1.5503,1.5503
20101229,204700,1.5503,1.5503,1.5502,1.5503
20101229,204800,1.5503,1.5503,1.5502,1.5502
20101229,204900,1.5502,1.5504,1.5501,1.5501
20101229,205000,1.55,1.5501,1.5499,1.5499
20101229,205100,1.55,1.5501,1.55,1.55
20101229,205200,1.5499,1.5499,1.5497,1.5498
20101229,205300,1.5498,1.5498,1.5497,1.5498
20101229,205400,1.5498,1.55,1.5498,1.5499
20101229,205500,1.55,1.55,1.5498,1.5498
20101229,205600,1.55,1.55,1.5498,1.5498
20101229,205700,1.55,1.5501,1.55,1.55
20101229,205800,1.5499,1.5499,1.5495,1.5495
20101229,205900,1.5495,1.5496,1.5495,1.5496
20101229,210000,1.5495,1.5496,1.5494,1.5495
20101229,210100,1.5495,1.5496,1.5495,1.5495
20101229,210200,1.5495,1.5495,1.5495,1.5495
20101229,210300,1.5495,1.5496,1.5495,1.5495
20101229,210400,1.5494,1.5495,1.5493,1.5493
20101229,210500,1.5494,1.5494,1.5493,1.5494
20101229,210600,1.5493,1.5493,1.5492,1.5492
20101229,210700,1.5493,1.5493,1.5491,1.5491
20101229,210800,1.549,1.5491,1.5488,1.5488
20101229,210900,1.5489,1.549,1.5488,1.5489
20101229,211000,1.5489,1.5489,1.5487,1.5487
20101229,211100,1.5488,1.5493,1.5488,1.5492
20101229,211200,1.5492,1.5492,1.5491,1.5491
20101229,211300,1.5491,1.5493,1.5489,1.5493
20101229,211400,1.5493,1.5494,1.5493,1.5494
20101229,211500,1.5493,1.5495,1.5493,1.5495
20101229,211600,1.5496,1.5498,1.5496,1.5498
20101229,211700,1.5497,1.5497,1.5497,1.5497
20101229,211800,1.5497,1.5497,1.5495,1.5495
20101229,211900,1.5496,1.5497,1.5496,1.5496
20101229,212000,1.5496,1.5496,1.5495,1.5496
20101229,212100,1.5496,1.5497,1.5496,1.5497
20101229,212200,1.5496,1.5497,1.5496,1.5497
20101229,212300,1.5497,1.5498,1.5497,1.5498
20101229,212400,1.5498,1.5499,1.5497,1.5499
20101229,212500,1.5499,1.5499,1.5497,1.5497
20101229,212600,1.5497,1.5498,1.5497,1.5498
20101229,212700,1.5499,1.5499,1.5498,1.5498
20101229,212800,1.5499,1.5499,1.5498,1.5498
20101229,212900,1.5498,1.5498,1.5498,1.5498
20101229,213000,1.5498,1.5498,1.5497,1.5497
20101229,213100,1.5497,1.5497,1.5497,1.5497
20101229,213200,1.5497,1.5498,1.5497,1.5498
20101229,213300,1.5497,1.5497,1.5497,1.5497
20101229,213400,1.5498,1.5498,1.5498,1.5498
20101229,213500,1.5498,1.5498,1.5498,1.5498
20101229,213600,1.5499,1.5499,1.5499,1.5499
20101229,213700,1.5499,1.5499,1.5499,1.5499
20101229,213800,1.5499,1.5499,1.5498,1.5498
20101229,213900,1.5498,1.5499,1.5496,1.5499
20101229,214000,1.5499,1.5499,1.5498,1.5498
20101229,214100,1.5498,1.5498,1.5493,1.5493
20101229,214200,1.5493,1.5493,1.5492,1.5493
20101229,214300,1.5493,1.5493,1.5493,1.5493
20101229,214400,1.5493,1.5493,1.5491,1.5493
20101229,214500,1.5493,1.5494,1.5493,1.5494
20101229,214600,1.5495,1.5496,1.5494,1.5495
20101229,214700,1.5495,1.5495,1.5493,1.5493
20101229,214800,1.5493,1.5495,1.5492,1.5495
20101229,214900,1.5496,1.5496,1.5495,1.5495
20101229,215000,1.5495,1.5495,1.5495,1.5495
20101229,215100,1.5495,1.5495,1.5494,1.5494
20101229,215200,1.5495,1.5495,1.5494,1.5494
20101229,215300,1.5494,1.5495,1.5494,1.5495
20101229,215400,1.5495,1.5495,1.5495,1.5495
20101229,215500,1.5496,1.5496,1.5495,1.5495
20101229,215600,1.5495,1.5495,1.5495,1.5495
20101229,215700,1.5496,1.5498,1.5496,1.5496
20101229,215800,1.5495,1.5496,1.5495,1.5496
20101229,215900,1.5495,1.5497,1.5495,1.5497
20101229,220000,1.5496,1.5498,1.5496,1.5498
20101229,220100,1.5498,1.5499,1.5498,1.5499
20101229,220200,1.5498,1.5498,1.5496,1.5497
20101229,220300,1.5496,1.5496,1.5496,1.5496
20101229,220400,1.5495,1.5497,1.5495,1.5497
20101229,220500,1.5497,1.5497,1.5495,1.5495
20101229,220600,1.5495,1.5496,1.5495,1.5496
20101229,220700,1.5496,1.5496,1.5496,1.5496
20101229,220800,1.5496,1.5497,1.5495,1.5495
20101229,220900,1.5496,1.5496,1.5496,1.5496
20101229,221000,1.5496,1.5497,1.5496,1.5497
20101229,221100,1.5497,1.5497,1.5495,1.5496
20101229,221200,1.5497,1.5498,1.5497,1.5497
20101229,221300,1.5495,1.5496,1.5495,1.5495
20101229,221400,1.5495,1.5495,1.5495,1.5495
20101229,221500,1.5495,1.5496,1.5495,1.5495
20101229,221600,1.5496,1.5504,1.5496,1.5504
20101229,221700,1.5504,1.5509,1.5504,1.5506
20101229,221800,1.5509,1.551,1.5501,1.5504
20101229,221900,1.5504,1.5504,1.5503,1.5503
20101229,222000,1.5502,1.5504,1.5502,1.5504
20101229,222100,1.5504,1.5504,1.5503,1.5503
20101229,222200,1.55,1.5501,1.55,1.5501
20101229,222300,1.5502,1.5503,1.5501,1.5503
20101229,222400,1.5503,1.5503,1.5502,1.5502
20101229,222500,1.5502,1.5502,1.5502,1.5502
20101229,222600,1.5502,1.5502,1.5502,1.5502
20101229,222700,1.5502,1.5503,1.5502,1.5503
20101229,222800,1.5504,1.5504,1.5502,1.5502
20101229,222900,1.5502,1.5502,1.5502,1.5502
20101229,223000,1.5502,1.5503,1.5501,1.5501
20101229,223100,1.55,1.55,1.5496,1.5496
20101229,223200,1.5497,1.5497,1.5497,1.5497
20101229,223300,1.5497,1.5497,1.5496,1.5497
20101229,223400,1.5498,1.5498,1.5497,1.5497
20101229,223500,1.5497,1.5497,1.5496,1.5496
20101229,223600,1.5496,1.5497,1.5495,1.5495
20101229,223700,1.5495,1.5495,1.5494,1.5494
20101229,223800,1.5494,1.5495,1.5494,1.5494
20101229,223900,1.5493,1.5493,1.5493,1.5493
20101229,224000,1.5495,1.5495,1.5494,1.5494
20101229,224100,1.5493,1.5493,1.5493,1.5493
20101229,224200,1.5494,1.5494,1.5494,1.5494
20101229,224300,1.5483,1.5483,1.5483,1.5483
20101229,224400,1.5485,1.5485,1.5485,1.5485
20101229,224600,1.5483,1.5483,1.5483,1.5483
20101229,224700,1.5492,1.5492,1.5492,1.5492
20101229,224800,1.5492,1.5492,1.5492,1.5492
20101229,224900,1.5492,1.5492,1.5492,1.5492
20101229,225000,1.5496,1.5496,1.5496,1.5496
20101229,225100,1.5498,1.5498,1.5498,1.5498
20101229,225300,1.5498,1.5499,1.5498,1.5499
20101229,225400,1.5498,1.5498,1.5498,1.5498
20101229,225600,1.5498,1.5498,1.5498,1.5498
20101229,225700,1.5498,1.5498,1.5497,1.5497
20101229,225800,1.5497,1.5498,1.5495,1.5495
20101229,225900,1.5496,1.5496,1.5496,1.5496
20101229,230000,1.5496,1.5496,1.5496,1.5496
20101229,230100,1.5496,1.5496,1.5496,1.5496
20101229,230300,1.5497,1.5497,1.5496,1.5496
20101229,230400,1.5495,1.5495,1.5495,1.5495
20101229,230500,1.5495,1.5495,1.5495,1.5495
20101229,230600,1.5496,1.5496,1.5496,1.5496
20101229,230800,1.5496,1.5496,1.5496,1.5496
20101229,230900,1.5495,1.5495,1.5495,1.5495
20101229,231100,1.5495,1.5495,1.5495,1.5495
20101229,231200,1.5496,1.5496,1.5496,1.5496
20101229,231400,1.5495,1.5495,1.5495,1.5495
20101229,231600,1.5495,1.5495,1.5495,1.5495
20101229,231700,1.5496,1.5496,1.5496,1.5496
20101229,231800,1.5496,1.5496,1.5496,1.5496
20101229,231900,1.5495,1.5495,1.5495,1.5495
20101229,232100,1.5495,1.5495,1.5495,1.5495
20101229,232300,1.5496,1.5496,1.5496,1.5496
20101229,232500,1.5497,1.5497,1.5496,1.5496
20101229,232600,1.5494,1.5494,1.5494,1.5494
20101229,232800,1.5494,1.5495,1.5494,1.5494
20101229,233000,1.5494,1.5494,1.5494,1.5494
20101229,233200,1.5494,1.5494,1.5494,1.5494
20101229,233300,1.5494,1.5494,1.5494,1.5494
20101229,233500,1.5494,1.5494,1.5494,1.5494
20101229,233600,1.5493,1.5494,1.5493,1.5494
20101229,233700,1.5494,1.5494,1.5492,1.5493
20101229,233800,1.5494,1.5495,1.5494,1.5495
20101229,233900,1.5494,1.5494,1.5494,1.5494
20101229,234100,1.5494,1.5494,1.5494,1.5494
20101229,234300,1.5494,1.5495,1.5494,1.5494
20101229,234400,1.5493,1.5493,1.5493,1.5493
20101229,234500,1.5497,1.5497,1.5497,1.5497
20101229,234700,1.5496,1.5496,1.5496,1.5496
20101229,234900,1.5495,1.5495,1.5495,1.5495
20101229,235000,1.5497,1.5497,1.5497,1.5497
20101229,235200,1.5498,1.5499,1.5498,1.5499
20101229,235300,1.55,1.55,1.55,1.55
20101229,235500,1.5498,1.5498,1.5498,1.5498
20101229,235700,1.5498,1.55,1.5497,1.5499
20101229,235800,1.5499,1.5499,1.5498,1.5498
20101229,235900,1.5498,1.5498,1.5498,1.5498
20101230,0,1.5498,1.55,1.5498,1.55
20101230,100,1.55,1.55,1.55,1.55
20101230,200,1.55,1.55,1.55,1.55
20101230,300,1.55,1.55,1.55,1.55
20101230,400,1.55,1.55,1.55,1.55
20101230,600,1.55,1.5501,1.55,1.5501
20101230,700,1.5497,1.5497,1.5497,1.5497
20101230,900,1.5498,1.5498,1.5497,1.5497
20101230,1000,1.55,1.55,1.55,1.55
20101230,1100,1.5503,1.5503,1.5503,1.5503
20101230,1200,1.5502,1.5502,1.5501,1.5502
20101230,1400,1.5504,1.5504,1.5504,1.5504
20101230,1600,1.5506,1.5506,1.5506,1.5506
20101230,1700,1.551,1.551,1.551,1.551
20101230,1900,1.5523,1.5523,1.5523,1.5523
20101230,2000,1.552,1.552,1.552,1.552
20101230,2100,1.552,1.552,1.552,1.552
20101230,2300,1.5517,1.5517,1.5517,1.5517
20101230,2500,1.5521,1.5521,1.5521,1.5521
20101230,2600,1.5521,1.5521,1.5521,1.5521
20101230,2800,1.552,1.5521,1.552,1.5521
20101230,2900,1.5522,1.5522,1.5522,1.5522
20101230,3100,1.5522,1.5522,1.5521,1.5522
20101230,3200,1.5522,1.5522,1.5522,1.5522
20101230,3300,1.552,1.552,1.552,1.552
20101230,3400,1.5518,1.5518,1.5518,1.5518
20101230,3500,1.552,1.552,1.552,1.552
20101230,3600,1.552,1.552,1.552,1.552
20101230,3800,1.552,1.552,1.552,1.552
20101230,3900,1.5518,1.5518,1.5518,1.5518
20101230,4000,1.5517,1.5517,1.5517,1.5517
20101230,4200,1.5517,1.5517,1.5514,1.5514
20101230,4300,1.5515,1.5516,1.5514,1.5515
20101230,4400,1.5519,1.5519,1.5519,1.5519
20101230,4500,1.552,1.552,1.552,1.552
20101230,4600,1.5519,1.5519,1.5519,1.5519
20101230,4800,1.5523,1.5523,1.5523,1.5523
20101230,4900,1.5523,1.5523,1.5523,1.5523
20101230,5000,1.5524,1.5524,1.5524,1.5524
20101230,5100,1.5525,1.5525,1.5525,1.5525
20101230,5200,1.5524,1.5524,1.5521,1.5524
20101230,5400,1.552,1.552,1.552,1.552
20101230,5500,1.552,1.552,1.552,1.552
20101230,5600,1.5519,1.5519,1.5519,1.5519
20101230,5700,1.5519,1.5519,1.5519,1.5519
20101230,5900,1.5518,1.5518,1.5516,1.5517
20101230,10000,1.5518,1.5518,1.5517,1.5518
20101230,10100,1.5518,1.5518,1.5518,1.5518
20101230,10300,1.5519,1.5519,1.5519,1.5519
20101230,10400,1.5524,1.5524,1.5524,1.5524
20101230,10500,1.5524,1.5524,1.5524,1.5524
20101230,10600,1.5524,1.5524,1.5524,1.5524
20101230,10700,1.5523,1.5523,1.5523,1.5523
20101230,10800,1.5523,1.5523,1.5523,1.5523
20101230,11000,1.5524,1.5524,1.5524,1.5524
20101230,11100,1.5525,1.5526,1.5525,1.5525
20101230,11200,1.5525,1.5525,1.5525,1.5525
20101230,11300,1.5525,1.5526,1.5525,1.5525
20101230,11400,1.5526,1.5526,1.5526,1.5526
20101230,11500,1.5526,1.5526,1.5526,1.5526
20101230,11700,1.5527,1.5527,1.5527,1.5527
20101230,11800,1.5525,1.5525,1.5525,1.5525
20101230,12000,1.5525,1.5525,1.5525,1.5525
20101230,12200,1.5525,1.5525,1.5525,1.5525
20101230,12300,1.5525,1.5526,1.5525,1.5526
20101230,12400,1.5526,1.5527,1.5526,1.5527
20101230,12500,1.5525,1.5527,1.5525,1.5525
20101230,12600,1.5525,1.5525,1.5524,1.5524
20101230,12700,1.5523,1.5523,1.5522,1.5522
20101230,12800,1.5522,1.5522,1.552,1.5521
20101230,12900,1.552,1.5522,1.552,1.5521
20101230,13000,1.5519,1.5519,1.5519,1.5519
20101230,13100,1.5519,1.5519,1.5519,1.5519
20101230,13300,1.5519,1.5519,1.5517,1.5517
20101230,13400,1.5518,1.552,1.5518,1.552
20101230,13500,1.552,1.5521,1.5519,1.5521
20101230,13600,1.552,1.552,1.5519,1.552
20101230,13700,1.5522,1.5522,1.5522,1.5522
20101230,13800,1.5523,1.5523,1.5523,1.5523
20101230,14000,1.5524,1.5524,1.5523,1.5523
20101230,14100,1.5524,1.5524,1.5523,1.5523
20101230,14200,1.5522,1.5522,1.5522,1.5522
20101230,14300,1.5522,1.5522,1.5522,1.5522
20101230,14400,1.552,1.552,1.552,1.552
20101230,14600,1.5519,1.5523,1.5519,1.5523
20101230,14700,1.5522,1.5522,1.5521,1.5521
20101230,14800,1.552,1.5522,1.552,1.5521
20101230,14900,1.5522,1.5522,1.5522,1.5522
20101230,15000,1.552,1.552,1.552,1.552
20101230,15200,1.552,1.552,1.552,1.552
20101230,15400,1.552,1.5521,1.5519,1.5521
20101230,15500,1.552,1.5521,1.552,1.552
20101230,15600,1.552,1.552,1.552,1.552
20101230,15700,1.552,1.5521,1.552,1.552
20101230,15800,1.5519,1.5519,1.5519,1.5519
20101230,15900,1.552,1.552,1.552,1.552
20101230,20000,1.5514,1.5514,1.5514,1.5514
20101230,20100,1.5515,1.5515,1.5515,1.5515
20101230,20300,1.5516,1.5516,1.5514,1.5516
20101230,20400,1.5517,1.5518,1.5515,1.5516
20101230,20500,1.5516,1.5516,1.5516,1.5516
20101230,20600,1.5515,1.5515,1.5515,1.5515
20101230,20700,1.5514,1.5514,1.5514,1.5514
20101230,20800,1.5515,1.5515,1.5515,1.5515
20101230,21000,1.5513,1.5513,1.5513,1.5513
20101230,21100,1.5514,1.5514,1.5514,1.5514
20101230,21300,1.5514,1.5514,1.5513,1.5513
20101230,21400,1.5512,1.5514,1.5512,1.5514
20101230,21600,1.5514,1.5515,1.5513,1.5515
20101230,21700,1.5514,1.5514,1.5514,1.5514
20101230,21800,1.5513,1.5513,1.5512,1.5513
20101230,22000,1.5513,1.5514,1.5513,1.5514
20101230,22100,1.5513,1.5513,1.5513,1.5513
20101230,22200,1.551,1.551,1.551,1.551
20101230,22400,1.5512,1.5512,1.5512,1.5512
20101230,22600,1.5512,1.5513,1.5512,1.5513
20101230,22700,1.5512,1.5512,1.5511,1.5512
20101230,22800,1.5513,1.5513,1.5513,1.5513
20101230,22900,1.5514,1.5514,1.5514,1.5514
20101230,23100,1.5513,1.5513,1.5513,1.5513
20101230,23300,1.5513,1.5513,1.5513,1.5513
20101230,23400,1.5511,1.5511,1.5511,1.5511
20101230,23500,1.5509,1.5509,1.5509,1.5509
20101230,23600,1.551,1.551,1.551,1.551
20101230,23800,1.5509,1.5509,1.5508,1.5509
20101230,23900,1.5508,1.5508,1.5508,1.5508
20101230,24100,1.5507,1.5507,1.5507,1.5507
20101230,24200,1.5507,1.5507,1.5507,1.5507
20101230,24300,1.5507,1.5507,1.5507,1.5507
20101230,24400,1.5508,1.5508,1.5508,1.5508
20101230,24500,1.5509,1.5509,1.5509,1.5509
20101230,24600,1.5511,1.5511,1.5511,1.5511
20101230,24800,1.5511,1.5511,1.551,1.551
20101230,24900,1.5511,1.5511,1.5509,1.551
20101230,25000,1.551,1.551,1.5509,1.5509
20101230,25100,1.5511,1.5511,1.5511,1.5511
20101230,25300,1.5511,1.5511,1.5509,1.5509
20101230,25400,1.551,1.551,1.551,1.551
20101230,25500,1.5509,1.551,1.5509,1.5509
20101230,25700,1.5509,1.551,1.5509,1.551
20101230,25800,1.5509,1.5509,1.5509,1.5509
20101230,30000,1.5509,1.551,1.5509,1.551
20101230,30100,1.551,1.551,1.5508,1.5509
20101230,30200,1.551,1.5511,1.551,1.551
20101230,30300,1.5511,1.5512,1.5509,1.5509
20101230,30400,1.5509,1.5511,1.5509,1.551
20101230,30500,1.551,1.5511,1.5509,1.5511
20101230,30600,1.5509,1.5509,1.5509,1.5509
20101230,30800,1.5508,1.551,1.5508,1.551
20101230,30900,1.5509,1.5509,1.5509,1.5509
20101230,31100,1.5508,1.5508,1.5508,1.5508
20101230,31300,1.5509,1.5509,1.5508,1.5508
20101230,31400,1.5508,1.5508,1.5507,1.5508
20101230,31500,1.5508,1.5508,1.5507,1.5508
20101230,31700,1.5507,1.5507,1.5507,1.5507
20101230,31800,1.5507,1.5507,1.5507,1.5507
20101230,32000,1.551,1.551,1.551,1.551
20101230,32100,1.551,1.551,1.551,1.551
20101230,32200,1.551,1.551,1.551,1.551
20101230,32300,1.5509,1.5509,1.5509,1.5509
20101230,32500,1.5509,1.5509,1.5509,1.5509
20101230,32600,1.5511,1.5511,1.5511,1.5511
20101230,32700,1.551,1.551,1.551,1.551
20101230,32900,1.5512,1.5512,1.5512,1.5512
20101230,33100,1.5512,1.5512,1.5512,1.5512
20101230,33200,1.5512,1.5512,1.5512,1.5512
20101230,33300,1.5512,1.5512,1.5512,1.5512
20101230,33500,1.551,1.5512,1.551,1.5511
20101230,33600,1.5512,1.5512,1.5512,1.5512
20101230,33700,1.551,1.551,1.551,1.551
20101230,33900,1.5512,1.5512,1.5512,1.5512
20101230,34100,1.5508,1.5508,1.5508,1.5508
20101230,34200,1.5508,1.5508,1.5508,1.5508
20101230,34400,1.5508,1.5508,1.5508,1.5508
20101230,34500,1.5508,1.5508,1.5508,1.5508
20101230,34600,1.5509,1.5509,1.5509,1.5509
20101230,34700,1.5509,1.5509,1.5509,1.5509
20101230,34900,1.5508,1.5509,1.5508,1.5509
20101230,35000,1.5509,1.5509,1.5508,1.5508
20101230,35100,1.5506,1.5506,1.5506,1.5506
20101230,35200,1.5506,1.5506,1.5506,1.5506
20101230,35400,1.5506,1.5506,1.5506,1.5506
20101230,35500,1.5504,1.5504,1.5504,1.5504
20101230,35600,1.5506,1.5506,1.5506,1.5506
20101230,35700,1.5506,1.5506,1.5506,1.5506
20101230,35800,1.5504,1.5504,1.5504,1.5504
20101230,35900,1.5504,1.5504,1.5504,1.5504
20101230,40000,1.5503,1.5503,1.5503,1.5503
20101230,40100,1.5504,1.5504,1.5504,1.5504
20101230,40200,1.5504,1.5504,1.5504,1.5504
20101230,40400,1.5504,1.5504,1.5504,1.5504
20101230,40600,1.5504,1.5504,1.5504,1.5504
20101230,40700,1.5504,1.5504,1.5504,1.5504
20101230,40800,1.5504,1.5504,1.5504,1.5504
20101230,41000,1.5506,1.5506,1.5504,1.5504
20101230,41100,1.5504,1.5504,1.5503,1.5503
20101230,41200,1.5503,1.5503,1.5503,1.5503
20101230,41400,1.5503,1.5503,1.5503,1.5503
20101230,41500,1.5502,1.5503,1.5502,1.5503
20101230,41600,1.5503,1.5504,1.5503,1.5504
20101230,41700,1.5503,1.5503,1.5502,1.5502
20101230,41800,1.5502,1.5502,1.5502,1.5502
20101230,41900,1.5503,1.5503,1.5503,1.5503
20101230,42000,1.5503,1.5504,1.5503,1.5503
20101230,42100,1.5504,1.5504,1.5504,1.5504
20101230,42300,1.5504,1.5504,1.5504,1.5504
20101230,42400,1.5504,1.5504,1.5504,1.5504
20101230,42600,1.5503,1.5504,1.5503,1.5504
20101230,42700,1.5502,1.5502,1.5502,1.5502
20101230,42900,1.5503,1.5503,1.5502,1.5503
20101230,43000,1.5503,1.5504,1.5503,1.5504
20101230,43100,1.5505,1.5505,1.5505,1.5505
20101230,43200,1.5506,1.5506,1.5506,1.5506
20101230,43300,1.5506,1.5506,1.5506,1.5506
20101230,43400,1.5506,1.5507,1.5506,1.5506
20101230,43600,1.5505,1.5505,1.5505,1.5505
20101230,43800,1.5504,1.5504,1.5504,1.5504
20101230,43900,1.5505,1.5505,1.5505,1.5505
20101230,44000,1.5506,1.5506,1.5506,1.5506
20101230,44200,1.5506,1.5506,1.5505,1.5506
20101230,44300,1.5506,1.5506,1.5506,1.5506
20101230,44400,1.5506,1.5507,1.5505,1.5506
20101230,44500,1.5506,1.5507,1.5506,1.5507
20101230,44600,1.5507,1.5507,1.5506,1.5506
20101230,44700,1.5507,1.5507,1.5507,1.5507
20101230,44800,1.5508,1.5508,1.5508,1.5508
20101230,45000,1.5507,1.5507,1.5507,1.5507
20101230,45200,1.5508,1.5508,1.5507,1.5507
20101230,45300,1.5507,1.5507,1.5507,1.5507
20101230,45400,1.5507,1.5508,1.5507,1.5507
20101230,45600,1.5508,1.5508,1.5508,1.5508
20101230,45700,1.5509,1.5509,1.5509,1.5509
20101230,45800,1.5509,1.5509,1.5509,1.5509
20101230,45900,1.5509,1.5509,1.5509,1.5509
20101230,50000,1.5509,1.5509,1.5509,1.5509
20101230,50100,1.5509,1.5509,1.5508,1.5509
20101230,50200,1.5508,1.5509,1.5508,1.5508
20101230,50300,1.5508,1.5508,1.5508,1.5508
20101230,50500,1.5506,1.5506,1.5506,1.5506
20101230,50700,1.5507,1.5507,1.5507,1.5507
20101230,50800,1.5507,1.5507,1.5507,1.5507
20101230,51000,1.5507,1.5508,1.5507,1.5507
20101230,51100,1.5508,1.5508,1.5508,1.5508
20101230,51200,1.5507,1.5508,1.5507,1.5508
20101230,51300,1.5508,1.5508,1.5507,1.5508
20101230,51400,1.5508,1.5508,1.5507,1.5507
20101230,51500,1.5507,1.5507,1.5507,1.5507
20101230,51600,1.5508,1.5508,1.5507,1.5507
20101230,51700,1.5507,1.551,1.5507,1.551
20101230,51800,1.551,1.551,1.5509,1.5509
20101230,51900,1.551,1.551,1.5508,1.5509
20101230,52000,1.5508,1.5509,1.5507,1.5507
20101230,52100,1.5506,1.5506,1.5506,1.5506
20101230,52300,1.5507,1.5507,1.5507,1.5507
20101230,52400,1.5506,1.551,1.5506,1.551
20101230,52500,1.5513,1.5513,1.5513,1.5513
20101230,52600,1.5513,1.5513,1.5512,1.5513
20101230,52700,1.5513,1.5513,1.5512,1.5513
20101230,52800,1.5511,1.5511,1.5511,1.5511
20101230,53000,1.5511,1.5511,1.5511,1.5511
20101230,53100,1.5511,1.5511,1.5511,1.5511
20101230,53300,1.5513,1.5513,1.5513,1.5513
20101230,53500,1.551,1.551,1.551,1.551
20101230,53600,1.551,1.551,1.551,1.551
20101230,53700,1.5509,1.5509,1.5509,1.5509
20101230,53800,1.5509,1.5509,1.5509,1.5509
20101230,54000,1.5511,1.5511,1.5511,1.5511
20101230,54200,1.551,1.551,1.5509,1.551
20101230,54300,1.5508,1.5508,1.5508,1.5508
20101230,54500,1.5508,1.551,1.5508,1.551
20101230,54600,1.5509,1.5511,1.5509,1.5511
20101230,54700,1.5513,1.5513,1.5513,1.5513
20101230,54800,1.551,1.551,1.551,1.551
20101230,55000,1.551,1.551,1.551,1.551
20101230,55100,1.551,1.551,1.551,1.551
20101230,55200,1.551,1.551,1.551,1.551
20101230,55400,1.5509,1.5509,1.5509,1.5509
20101230,55500,1.5511,1.5511,1.5511,1.5511
20101230,55600,1.551,1.551,1.551,1.551
20101230,55800,1.551,1.5511,1.551,1.5511
20101230,55900,1.5511,1.5511,1.551,1.5511
20101230,60000,1.551,1.5513,1.551,1.5513
20101230,60100,1.5512,1.5513,1.5511,1.5513
20101230,60200,1.5513,1.5513,1.5512,1.5512
20101230,60300,1.5512,1.5512,1.5512,1.5512
20101230,60400,1.5515,1.5515,1.5515,1.5515
20101230,60500,1.5515,1.5515,1.5515,1.5515
20101230,60700,1.5515,1.5515,1.5514,1.5515
20101230,60800,1.5515,1.5515,1.5515,1.5515
20101230,61000,1.5516,1.5517,1.5516,1.5517
20101230,61100,1.5517,1.5517,1.5517,1.5517
20101230,61200,1.5518,1.5518,1.5518,1.5518
20101230,61400,1.5516,1.5516,1.5516,1.5516
20101230,61600,1.5516,1.5516,1.5516,1.5516
20101230,61800,1.5517,1.5517,1.5517,1.5517
20101230,62000,1.5516,1.5517,1.5516,1.5517
20101230,62100,1.5517,1.5517,1.5517,1.5517
20101230,62200,1.5517,1.5517,1.5517,1.5517
20101230,62300,1.5517,1.5517,1.5516,1.5516
20101230,62400,1.5518,1.5518,1.5518,1.5518
20101230,62600,1.5517,1.5517,1.5517,1.5517
20101230,62700,1.5518,1.5518,1.5518,1.5518
20101230,62900,1.5519,1.5519,1.5519,1.5519
20101230,63000,1.5517,1.5517,1.5517,1.5517
20101230,63100,1.5517,1.5517,1.5517,1.5517
20101230,63200,1.5513,1.5513,1.5513,1.5513
20101230,63300,1.5514,1.5514,1.5514,1.5514
20101230,63400,1.5513,1.5513,1.5513,1.5513
20101230,63600,1.5514,1.5514,1.5514,1.5514
20101230,63700,1.5515,1.5515,1.5515,1.5515
20101230,63900,1.5516,1.5516,1.5516,1.5516
20101230,64100,1.5516,1.5516,1.5514,1.5515
20101230,64200,1.5515,1.5516,1.5515,1.5515
20101230,64300,1.5514,1.5516,1.5514,1.5516
20101230,64400,1.5515,1.5515,1.5515,1.5515
20101230,64500,1.5516,1.5516,1.5516,1.5516
20101230,64600,1.5513,1.5513,1.5513,1.5513
20101230,64700,1.5511,1.5511,1.5511,1.5511
20101230,64800,1.5512,1.5512,1.5512,1.5512
20101230,65000,1.5511,1.5511,1.5511,1.5511
20101230,65100,1.5511,1.5511,1.551,1.551
20101230,65200,1.5509,1.551,1.5508,1.551
20101230,65300,1.5509,1.5509,1.5508,1.5509
20101230,65400,1.5509,1.5509,1.5508,1.5509
20101230,65500,1.5507,1.5507,1.5507,1.5507
20101230,65700,1.5508,1.5508,1.5508,1.5508
20101230,65800,1.5508,1.5508,1.5508,1.5508
20101230,65900,1.5508,1.5508,1.5508,1.5508
20101230,70000,1.5507,1.5507,1.5507,1.5507
20101230,70100,1.5508,1.5508,1.5508,1.5508
20101230,70300,1.5512,1.5512,1.5512,1.5512
20101230,70400,1.5515,1.5515,1.5515,1.5515
20101230,70500,1.5516,1.5516,1.5516,1.5516
20101230,70600,1.5517,1.5517,1.5517,1.5517
20101230,70700,1.5517,1.5517,1.5517,1.5517
20101230,70900,1.5516,1.552,1.5515,1.5519
20101230,71100,1.5518,1.5518,1.5517,1.5517
20101230,71200,1.5517,1.5517,1.5516,1.5517
20101230,71300,1.5519,1.5519,1.5519,1.5519
20101230,71500,1.552,1.5521,1.5519,1.5521
20101230,71600,1.5525,1.5525,1.5525,1.5525
20101230,71700,1.5527,1.5527,1.5527,1.5527
20101230,71800,1.5531,1.5531,1.5531,1.5531
20101230,71900,1.5533,1.5533,1.5533,1.5533
20101230,72100,1.5529,1.5529,1.5529,1.5529
20101230,72300,1.5525,1.5525,1.5525,1.5525
20101230,72500,1.5524,1.5524,1.5522,1.5522
20101230,72600,1.5525,1.5525,1.5525,1.5525
20101230,72700,1.5525,1.5525,1.5525,1.5525
20101230,72900,1.5525,1.5526,1.5525,1.5526
20101230,73000,1.5527,1.5528,1.5527,1.5528
20101230,73100,1.5528,1.5528,1.5528,1.5528
20101230,73200,1.5526,1.5526,1.5526,1.5526
20101230,73300,1.5525,1.5525,1.5525,1.5525
20101230,73400,1.5524,1.5524,1.5524,1.5524
20101230,73600,1.5523,1.5525,1.5522,1.5524
20101230,73800,1.5524,1.5524,1.5524,1.5524
20101230,74000,1.5519,1.5519,1.5519,1.5519
20101230,74100,1.5518,1.5518,1.5518,1.5518
20101230,74200,1.5519,1.5519,1.5519,1.5519
20101230,74300,1.552,1.5521,1.552,1.5521
20101230,74400,1.5521,1.5521,1.5521,1.5521
20101230,74500,1.5523,1.5523,1.5523,1.5523
20101230,74700,1.5522,1.5522,1.552,1.552
20101230,74800,1.552,1.5521,1.5519,1.5519
20101230,74900,1.5518,1.5519,1.5517,1.5519
20101230,75000,1.5518,1.5519,1.5518,1.5518
20101230,75100,1.5518,1.5519,1.5518,1.5518
20101230,75200,1.5518,1.5518,1.5518,1.5518
20101230,75300,1.5518,1.5518,1.5518,1.5518
20101230,75400,1.5517,1.5517,1.5517,1.5517
20101230,75500,1.5518,1.5518,1.5518,1.5518
20101230,75700,1.5519,1.5519,1.5517,1.5518
20101230,75800,1.5514,1.5514,1.5514,1.5514
20101230,75900,1.551,1.551,1.551,1.551
20101230,80000,1.5507,1.5507,1.5507,1.5507
20101230,80100,1.5517,1.5517,1.5517,1.5517
20101230,80200,1.5517,1.5517,1.5517,1.5517
20101230,80300,1.5515,1.5515,1.5515,1.5515
20101230,80400,1.5518,1.5518,1.5518,1.5518
20101230,80500,1.5516,1.5516,1.5516,1.5516
20101230,80600,1.5511,1.5511,1.5511,1.5511
20101230,80700,1.5511,1.5511,1.5511,1.5511
20101230,80800,1.5518,1.5518,1.5518,1.5518
20101230,80900,1.5517,1.5517,1.5517,1.5517
20101230,81000,1.5515,1.5515,1.5515,1.5515
20101230,81100,1.5514,1.5514,1.5514,1.5514
20101230,81200,1.5516,1.5516,1.5516,1.5516
20101230,81400,1.5514,1.5514,1.5514,1.5514
20101230,81500,1.5514,1.5514,1.5514,1.5514
20101230,81700,1.5513,1.5513,1.5512,1.5513
20101230,81800,1.5511,1.5511,1.5511,1.5511
20101230,81900,1.5511,1.5511,1.5511,1.5511
20101230,82000,1.551,1.551,1.551,1.551
20101230,82100,1.5511,1.5511,1.5511,1.5511
20101230,82200,1.5509,1.5509,1.5509,1.5509
20101230,82300,1.5508,1.5509,1.5508,1.5508
20101230,82400,1.5507,1.5507,1.5507,1.5507
20101230,82500,1.5503,1.5503,1.5503,1.5503
20101230,82600,1.5504,1.5504,1.5504,1.5504
20101230,82800,1.5502,1.5502,1.5502,1.5502
20101230,82900,1.55,1.55,1.55,1.55
20101230,83000,1.5501,1.5501,1.5501,1.5501
20101230,83100,1.5502,1.5502,1.5502,1.5502
20101230,83200,1.5501,1.5505,1.5501,1.5502
20101230,83300,1.55,1.55,1.55,1.55
20101230,83500,1.55,1.55,1.5499,1.55
20101230,83600,1.5504,1.5504,1.5504,1.5504
20101230,83700,1.5506,1.5506,1.5506,1.5506
20101230,83900,1.5506,1.5506,1.5506,1.5506
20101230,84100,1.5507,1.5507,1.5506,1.5506
20101230,84200,1.5505,1.5506,1.5504,1.5504
20101230,84300,1.5505,1.5505,1.5504,1.5505
20101230,84400,1.5504,1.5504,1.5503,1.5504
20101230,84500,1.5505,1.5505,1.5501,1.5501
20101230,84600,1.5501,1.5501,1.5501,1.5501
20101230,84800,1.5498,1.5498,1.5498,1.5498
20101230,84900,1.5495,1.5495,1.5495,1.5495
20101230,85100,1.5486,1.5486,1.5486,1.5486
20101230,85300,1.5489,1.5489,1.5489,1.5489
20101230,85400,1.5488,1.5488,1.5488,1.5488
20101230,85600,1.5485,1.5485,1.5485,1.5485
20101230,85700,1.5487,1.5487,1.5487,1.5487
20101230,85800,1.5488,1.5495,1.5488,1.5488
20101230,85900,1.5496,1.5496,1.5496,1.5496
20101230,90000,1.5496,1.5496,1.5496,1.5496
20101230,90100,1.5494,1.5494,1.5494,1.5494
20101230,90300,1.5494,1.5494,1.5494,1.5494
20101230,90500,1.5494,1.5494,1.5494,1.5494
20101230,90600,1.5495,1.5496,1.5495,1.5495
20101230,90700,1.5496,1.5496,1.5496,1.5496
20101230,90800,1.5495,1.5495,1.5495,1.5495
20101230,91000,1.549,1.549,1.549,1.549
20101230,91200,1.5494,1.5494,1.5494,1.5494
20101230,91400,1.5493,1.5493,1.5493,1.5493
20101230,91600,1.5495,1.5495,1.5495,1.5495
20101230,91800,1.5495,1.5495,1.5495,1.5495
20101230,91900,1.5497,1.5497,1.5497,1.5497
20101230,92000,1.5494,1.5494,1.5494,1.5494
20101230,92200,1.5492,1.5492,1.5492,1.5492
20101230,92300,1.549,1.549,1.549,1.549
20101230,92400,1.5492,1.5492,1.5492,1.5492
20101230,92500,1.5492,1.5492,1.5492,1.5492
20101230,92600,1.5488,1.5488,1.5488,1.5488
20101230,92700,1.5488,1.5488,1.5488,1.5488
20101230,92800,1.5493,1.5493,1.5493,1.5493
20101230,92900,1.5493,1.5493,1.5493,1.5493
20101230,93100,1.549,1.549,1.549,1.549
20101230,93200,1.5489,1.5489,1.5489,1.5489
20101230,93400,1.5487,1.549,1.5487,1.549
20101230,93500,1.5487,1.5487,1.5487,1.5487
20101230,93700,1.5485,1.5485,1.5485,1.5485
20101230,93800,1.5486,1.5486,1.5486,1.5486
20101230,93900,1.5489,1.5489,1.5489,1.5489
20101230,94000,1.5488,1.5488,1.5488,1.5488
20101230,94100,1.5488,1.549,1.5488,1.5488
20101230,94300,1.549,1.5495,1.549,1.5495
20101230,94400,1.5493,1.5493,1.5493,1.5493
20101230,94600,1.5506,1.5506,1.5506,1.5506
20101230,94700,1.5504,1.5504,1.5504,1.5504
20101230,94900,1.5504,1.5504,1.5504,1.5504
20101230,95000,1.5504,1.5504,1.5504,1.5504
20101230,95200,1.5504,1.5504,1.5503,1.5503
20101230,95300,1.5502,1.5502,1.5502,1.5502
20101230,95500,1.5504,1.5504,1.5504,1.5504
20101230,95700,1.5505,1.5505,1.5505,1.5505
20101230,95800,1.5504,1.5504,1.5504,1.5504
20101230,100000,1.5502,1.5502,1.5502,1.5502
20101230,100200,1.5501,1.5501,1.5501,1.5501
20101230,100300,1.5502,1.5502,1.5502,1.5502
20101230,100400,1.5501,1.5501,1.5501,1.5501
20101230,100600,1.5501,1.5502,1.5501,1.5502
20101230,100700,1.5501,1.5501,1.5501,1.5501
20101230,100900,1.55,1.5502,1.55,1.5502
20101230,101000,1.5501,1.5502,1.55,1.5501
20101230,101100,1.5501,1.5502,1.5501,1.5501
20101230,101200,1.5498,1.5498,1.5498,1.5498
20101230,101300,1.5497,1.5497,1.5497,1.5497
20101230,101400,1.5495,1.5495,1.5495,1.5495
20101230,101500,1.5494,1.5494,1.5494,1.5494
20101230,101700,1.5494,1.5494,1.5494,1.5494
20101230,101800,1.5494,1.5494,1.549,1.549
20101230,101900,1.5498,1.5498,1.5498,1.5498
20101230,102100,1.5497,1.5497,1.5497,1.5497
20101230,102200,1.5498,1.5498,1.5498,1.5498
20101230,102400,1.5488,1.5488,1.5488,1.5488
20101230,102600,1.5487,1.5487,1.548,1.5482
20101230,102700,1.5462,1.5462,1.5462,1.5462
20101230,102800,1.546,1.546,1.546,1.546
20101230,102900,1.5466,1.5466,1.5466,1.5466
20101230,103000,1.5466,1.5466,1.5466,1.5466
20101230,103100,1.5459,1.5459,1.5459,1.5459
20101230,103200,1.5459,1.5459,1.5459,1.5459
20101230,103300,1.5459,1.5459,1.5459,1.5459
20101230,103400,1.5461,1.5461,1.5461,1.5461
20101230,103500,1.5465,1.5465,1.5465,1.5465
20101230,103600,1.5469,1.5469,1.5469,1.5469
20101230,103700,1.5469,1.5469,1.5469,1.5469
20101230,103900,1.5468,1.5471,1.5468,1.5468
20101230,104000,1.5469,1.5469,1.5465,1.5465
20101230,104100,1.5462,1.5462,1.5462,1.5462
20101230,104300,1.5463,1.5464,1.546,1.5462
20101230,104400,1.5455,1.5455,1.5455,1.5455
20101230,104500,1.5453,1.5453,1.5453,1.5453
20101230,104600,1.5452,1.5452,1.5452,1.5452
20101230,104700,1.5451,1.5451,1.5451,1.5451
20101230,104900,1.5451,1.5451,1.5451,1.5451
20101230,105000,1.5452,1.5452,1.5452,1.5452
20101230,105100,1.5451,1.5451,1.5451,1.5451
20101230,105200,1.5449,1.5449,1.5449,1.5449
20101230,105300,1.5449,1.5449,1.5449,1.5449
20101230,105500,1.5448,1.5448,1.5448,1.5448
20101230,105600,1.545,1.545,1.545,1.545
20101230,105800,1.5451,1.5451,1.545,1.545
20101230,105900,1.545,1.545,1.545,1.545
20101230,110000,1.5449,1.5449,1.5449,1.5449
20101230,110200,1.545,1.545,1.5445,1.5445
20101230,110300,1.5445,1.5445,1.5443,1.5444
20101230,110400,1.5444,1.5444,1.5444,1.5444
20101230,110500,1.5439,1.5439,1.5439,1.5439
20101230,110700,1.544,1.5442,1.544,1.5441
20101230,110800,1.5442,1.5442,1.5434,1.5435
20101230,110900,1.5434,1.5434,1.5434,1.5434
20101230,111100,1.5435,1.5435,1.5435,1.5435
20101230,111300,1.5434,1.5435,1.5431,1.5432
20101230,111400,1.5429,1.5429,1.5429,1.5429
20101230,111500,1.5427,1.5427,1.5427,1.5427
20101230,111700,1.5424,1.5424,1.5424,1.5424
20101230,111800,1.5424,1.5425,1.5424,1.5424
20101230,112000,1.5425,1.5425,1.5423,1.5423
20101230,112100,1.5424,1.5427,1.5424,1.5427
20101230,112200,1.5426,1.5426,1.5426,1.5426
20101230,112300,1.542,1.542,1.542,1.542
20101230,112400,1.5415,1.5415,1.5415,1.5415
20101230,112500,1.5413,1.5413,1.5413,1.5413
20101230,112600,1.5415,1.5415,1.5415,1.5415
20101230,112800,1.5421,1.5421,1.5421,1.5421
20101230,112900,1.5422,1.5422,1.5422,1.5422
20101230,113000,1.5423,1.5423,1.5423,1.5423
20101230,113100,1.5424,1.5424,1.5424,1.5424
20101230,113200,1.5424,1.5424,1.5424,1.5424
20101230,113300,1.5422,1.5422,1.5422,1.5422
20101230,113400,1.5424,1.5424,1.5424,1.5424
20101230,113600,1.5423,1.5424,1.5422,1.5424
20101230,113700,1.5423,1.5423,1.5423,1.5423
20101230,113800,1.5429,1.5429,1.5429,1.5429
20101230,114000,1.5428,1.5431,1.5427,1.5428
20101230,114100,1.5424,1.5424,1.5424,1.5424
20101230,114300,1.5426,1.5426,1.5426,1.5426
20101230,114400,1.5426,1.5426,1.5426,1.5426
20101230,114500,1.5426,1.5426,1.5426,1.5426
20101230,114600,1.5427,1.5428,1.5427,1.5427
20101230,114700,1.5428,1.5428,1.5428,1.5428
20101230,114800,1.5425,1.5425,1.5425,1.5425
20101230,114900,1.5421,1.5421,1.5421,1.5421
20101230,115100,1.5421,1.5421,1.5421,1.5421
20101230,115200,1.5425,1.5425,1.5425,1.5425
20101230,115300,1.5425,1.5425,1.5425,1.5425
20101230,115400,1.5424,1.5424,1.5424,1.5424
20101230,115500,1.5422,1.5422,1.5422,1.5422
20101230,115700,1.5423,1.5423,1.5423,1.5423
20101230,115800,1.5427,1.5427,1.5427,1.5427
20101230,115900,1.5432,1.5432,1.5432,1.5432
20101230,120000,1.543,1.543,1.543,1.543
20101230,120100,1.5433,1.5433,1.5433,1.5433
20101230,120200,1.5436,1.5436,1.5436,1.5436
20101230,120300,1.5437,1.5437,1.5437,1.5437
20101230,120400,1.5438,1.5443,1.5438,1.5438
20101230,120500,1.5441,1.5441,1.5441,1.5441
20101230,120700,1.5443,1.5443,1.5443,1.5443
20101230,120900,1.5442,1.5443,1.5441,1.5442
20101230,121000,1.5444,1.5444,1.5444,1.5444
20101230,121100,1.5442,1.5442,1.5442,1.5442
20101230,121200,1.5441,1.5441,1.5441,1.5441
20101230,121300,1.5436,1.5436,1.5436,1.5436
20101230,121400,1.5433,1.5433,1.5433,1.5433
20101230,121500,1.5428,1.5428,1.5428,1.5428
20101230,121700,1.5428,1.543,1.5428,1.5428
20101230,121800,1.5429,1.543,1.5429,1.5429
20101230,122000,1.543,1.5438,1.5429,1.5438
20101230,122100,1.5436,1.5436,1.5436,1.5436
20101230,122300,1.5437,1.5437,1.5436,1.5436
20101230,122400,1.5435,1.5436,1.5435,1.5435
20101230,122500,1.5436,1.5436,1.5435,1.5436
20101230,122600,1.5434,1.5434,1.5434,1.5434
20101230,122700,1.5432,1.5432,1.5432,1.5432
20101230,122800,1.5433,1.5433,1.5433,1.5433
20101230,123000,1.5433,1.5433,1.5433,1.5433
20101230,123100,1.5435,1.5435,1.5435,1.5435
20101230,123200,1.5437,1.5437,1.5437,1.5437
20101230,123400,1.5441,1.5441,1.5441,1.5441
20101230,123600,1.5441,1.5445,1.5436,1.5443
20101230,123800,1.5432,1.5432,1.5432,1.5432
20101230,124000,1.5433,1.5438,1.5432,1.5438
20101230,124100,1.5438,1.5438,1.5438,1.5438
20101230,124300,1.5444,1.5444,1.5444,1.5444
20101230,124400,1.5441,1.5441,1.5441,1.5441
20101230,124600,1.5443,1.5443,1.5443,1.5443
20101230,124800,1.5438,1.5438,1.5438,1.5438
20101230,125000,1.5438,1.544,1.5438,1.544
20101230,125100,1.5439,1.544,1.5438,1.5439
20101230,125200,1.5438,1.5438,1.5438,1.5438
20101230,125300,1.5436,1.5436,1.5436,1.5436
20101230,125500,1.5435,1.5435,1.5435,1.5435
20101230,125700,1.5434,1.5434,1.5433,1.5433
20101230,125800,1.5433,1.5433,1.5433,1.5433
20101230,125900,1.5427,1.5427,1.5427,1.5427
20101230,130000,1.543,1.543,1.543,1.543
20101230,130100,1.5431,1.5431,1.5431,1.5431
20101230,130200,1.5436,1.5436,1.5436,1.5436
20101230,130400,1.5436,1.544,1.5436,1.544
20101230,130500,1.544,1.544,1.5438,1.5438
20101230,130600,1.5439,1.5442,1.5439,1.544
20101230,130700,1.5447,1.5447,1.5447,1.5447
20101230,130800,1.5446,1.5446,1.5446,1.5446
20101230,131000,1.5446,1.5446,1.5446,1.5446
20101230,131200,1.5442,1.5442,1.5442,1.5442
20101230,131300,1.5442,1.5442,1.5442,1.5442
20101230,131400,1.5438,1.5438,1.5438,1.5438
20101230,131500,1.5434,1.5434,1.5434,1.5434
20101230,131600,1.5434,1.5434,1.5434,1.5434
20101230,131800,1.5433,1.5433,1.5432,1.5432
20101230,131900,1.5433,1.5433,1.5433,1.5433
20101230,132000,1.5428,1.5428,1.5428,1.5428
20101230,132200,1.5427,1.5427,1.5422,1.5425
20101230,132300,1.5426,1.5429,1.5426,1.5428
20101230,132400,1.5421,1.5421,1.5421,1.5421
20101230,132600,1.5415,1.5415,1.5415,1.5415
20101230,132700,1.5412,1.5412,1.5412,1.5412
20101230,132800,1.5415,1.5415,1.5415,1.5415
20101230,132900,1.5416,1.5416,1.5416,1.5416
20101230,133000,1.5404,1.5404,1.5404,1.5404
20101230,133100,1.5409,1.5409,1.5409,1.5409
20101230,133200,1.5415,1.5415,1.5415,1.5415
20101230,133300,1.5419,1.5419,1.5419,1.5419
20101230,133400,1.542,1.542,1.542,1.542
20101230,133500,1.5424,1.5424,1.5424,1.5424
20101230,133700,1.5428,1.5428,1.5428,1.5428
20101230,133800,1.5426,1.5426,1.5426,1.5426
20101230,133900,1.5426,1.5426,1.5426,1.5426
20101230,134000,1.5424,1.5424,1.5424,1.5424
20101230,134200,1.5422,1.5422,1.5422,1.5422
20101230,134300,1.5416,1.5416,1.5416,1.5416
20101230,134500,1.5416,1.5416,1.5411,1.5411
20101230,134600,1.5405,1.5405,1.5405,1.5405
20101230,134700,1.5402,1.5402,1.5402,1.5402
20101230,134800,1.5401,1.5401,1.5401,1.5401
20101230,135000,1.5402,1.5402,1.5402,1.5402
20101230,135100,1.5402,1.5402,1.5402,1.5402
20101230,135300,1.5401,1.5401,1.5401,1.5401
20101230,135400,1.5404,1.5404,1.5404,1.5404
20101230,135500,1.5407,1.5407,1.5407,1.5407
20101230,135700,1.5415,1.5415,1.5415,1.5415
20101230,135800,1.5412,1.5412,1.5412,1.5412
20101230,135900,1.5417,1.5417,1.5417,1.5417
20101230,140000,1.5426,1.5426,1.5426,1.5426
20101230,140100,1.5425,1.5425,1.5425,1.5425
20101230,140200,1.5425,1.5425,1.5425,1.5425
20101230,140300,1.5424,1.5424,1.5424,1.5424
20101230,140400,1.5421,1.5421,1.5421,1.5421
20101230,140500,1.5419,1.5419,1.5419,1.5419
20101230,140700,1.5424,1.5424,1.5424,1.5424
20101230,140800,1.5423,1.5423,1.5423,1.5423
20101230,140900,1.5416,1.5416,1.5416,1.5416
20101230,141000,1.5417,1.5417,1.5417,1.5417
20101230,141100,1.5418,1.5419,1.5418,1.5418
20101230,141200,1.5417,1.5417,1.5417,1.5417
20101230,141300,1.5418,1.5418,1.5418,1.5418
20101230,141400,1.542,1.542,1.542,1.542
20101230,141500,1.5423,1.5423,1.5423,1.5423
20101230,141600,1.5419,1.5419,1.5419,1.5419
20101230,141800,1.542,1.5423,1.542,1.5423
20101230,141900,1.5419,1.5419,1.5419,1.5419
20101230,142000,1.5418,1.5418,1.5418,1.5418
20101230,142100,1.5421,1.5421,1.5421,1.5421
20101230,142200,1.5422,1.5422,1.5422,1.5422
20101230,142300,1.5422,1.5424,1.5422,1.5422
20101230,142400,1.5423,1.5423,1.5423,1.5423
20101230,142500,1.5419,1.5419,1.5419,1.5419
20101230,142600,1.5419,1.5422,1.5419,1.5419
20101230,142700,1.5422,1.5422,1.5422,1.5422
20101230,142900,1.5421,1.5421,1.5419,1.542
20101230,143100,1.5418,1.5418,1.5418,1.5418
20101230,143200,1.5419,1.5419,1.5419,1.5419
20101230,143300,1.5421,1.5421,1.5421,1.5421
20101230,143400,1.5422,1.5422,1.5422,1.5422
20101230,143600,1.5424,1.5424,1.5424,1.5424
20101230,143700,1.5424,1.5424,1.5424,1.5424
20101230,143800,1.5423,1.5423,1.5423,1.5423
20101230,144000,1.5422,1.5423,1.542,1.542
20101230,144200,1.5424,1.5424,1.5424,1.5424
20101230,144300,1.5425,1.5425,1.5425,1.5425
20101230,144400,1.5427,1.5427,1.5427,1.5427
20101230,144500,1.5422,1.5422,1.5422,1.5422
20101230,144600,1.5426,1.5426,1.5426,1.5426
20101230,144700,1.5426,1.5426,1.5426,1.5426
20101230,144800,1.5424,1.5424,1.5424,1.5424
20101230,144900,1.5429,1.5429,1.5429,1.5429
20101230,145000,1.5429,1.5429,1.5429,1.5429
20101230,145100,1.5434,1.5434,1.5434,1.5434
20101230,145200,1.5435,1.5435,1.5435,1.5435
20101230,145400,1.5439,1.5439,1.5439,1.5439
20101230,145500,1.5441,1.5441,1.5441,1.5441
20101230,145600,1.5445,1.5445,1.5445,1.5445
20101230,145700,1.5461,1.5461,1.5461,1.5461
20101230,145800,1.5459,1.5459,1.5459,1.5459
20101230,145900,1.546,1.546,1.546,1.546
20101230,150000,1.546,1.546,1.546,1.546
20101230,150100,1.5456,1.5456,1.5456,1.5456
20101230,150200,1.5457,1.5457,1.5457,1.5457
20101230,150300,1.5452,1.5452,1.5452,1.5452
20101230,150500,1.5449,1.5449,1.5449,1.5449
20101230,150600,1.5445,1.5445,1.5445,1.5445
20101230,150700,1.5445,1.5445,1.5445,1.5445
20101230,150900,1.5445,1.5446,1.5442,1.5444
20101230,151000,1.5445,1.5445,1.5445,1.5445
20101230,151200,1.5444,1.5444,1.5444,1.5444
20101230,151300,1.5442,1.5442,1.5442,1.5442
20101230,151500,1.5443,1.5443,1.5441,1.5442
20101230,151600,1.5443,1.5445,1.5443,1.5443
20101230,151700,1.5444,1.5446,1.5443,1.5443
20101230,151800,1.5443,1.5443,1.5443,1.5443
20101230,152000,1.5438,1.5438,1.5438,1.5438
20101230,152200,1.5438,1.5438,1.5438,1.5438
20101230,152300,1.5432,1.5432,1.5432,1.5432
20101230,152400,1.5431,1.5431,1.5431,1.5431
20101230,152500,1.5433,1.5433,1.5433,1.5433
20101230,152600,1.5434,1.5434,1.5434,1.5434
20101230,152700,1.5432,1.5432,1.5432,1.5432
20101230,152800,1.5431,1.5431,1.5431,1.5431
20101230,152900,1.543,1.543,1.5427,1.543
20101230,153100,1.5416,1.5416,1.5416,1.5416
20101230,153200,1.541,1.541,1.541,1.541
20101230,153300,1.5408,1.5408,1.5408,1.5408
20101230,153500,1.5405,1.5405,1.5405,1.5405
20101230,153600,1.5408,1.5408,1.5408,1.5408
20101230,153800,1.54,1.54,1.54,1.54
20101230,153900,1.5396,1.5396,1.5396,1.5396
20101230,154100,1.5397,1.5397,1.5396,1.5397
20101230,154200,1.5394,1.5394,1.5394,1.5394
20101230,154400,1.5394,1.5394,1.5394,1.5394
20101230,154500,1.5402,1.5402,1.5402,1.5402
20101230,154700,1.5402,1.5402,1.5402,1.5402
20101230,154800,1.5406,1.5406,1.5406,1.5406
20101230,154900,1.5405,1.5405,1.5403,1.5405
20101230,155000,1.5402,1.5402,1.5402,1.5402
20101230,155200,1.5405,1.5405,1.5405,1.5405
20101230,155300,1.5403,1.5403,1.5403,1.5403
20101230,155400,1.5404,1.5404,1.5404,1.5404
20101230,155500,1.5395,1.5395,1.5395,1.5395
20101230,155600,1.5394,1.5394,1.5394,1.5394
20101230,155700,1.5392,1.5392,1.5392,1.5392
20101230,155800,1.5388,1.5388,1.5388,1.5388
20101230,160000,1.5394,1.5394,1.5394,1.5394
20101230,160100,1.5396,1.5396,1.5396,1.5396
20101230,160300,1.5396,1.5399,1.5395,1.5395
20101230,160500,1.5398,1.5398,1.5398,1.5398
20101230,160600,1.5392,1.5392,1.5392,1.5392
20101230,160700,1.5391,1.5391,1.5391,1.5391
20101230,160800,1.5388,1.5388,1.5388,1.5388
20101230,161000,1.5384,1.5384,1.5384,1.5384
20101230,161200,1.5385,1.5385,1.5385,1.5385
20101230,161300,1.5384,1.5384,1.5383,1.5384
20101230,161400,1.5386,1.5386,1.5386,1.5386
20101230,161500,1.5388,1.5388,1.5388,1.5388
20101230,161600,1.5384,1.5384,1.5384,1.5384
20101230,161700,1.5383,1.5383,1.5383,1.5383
20101230,161900,1.5381,1.5381,1.5381,1.5381
20101230,162000,1.5376,1.5376,1.5376,1.5376
20101230,162100,1.5375,1.5375,1.5375,1.5375
20101230,162200,1.5381,1.5381,1.5381,1.5381
20101230,162300,1.5376,1.5376,1.5376,1.5376
20101230,162400,1.5375,1.5375,1.5375,1.5375
20101230,162600,1.5386,1.5386,1.5386,1.5386
20101230,162700,1.5382,1.5382,1.5382,1.5382
20101230,162800,1.5382,1.5382,1.5382,1.5382
20101230,162900,1.5384,1.5384,1.5384,1.5384
20101230,163000,1.5387,1.5387,1.5387,1.5387
20101230,163200,1.5386,1.5393,1.5386,1.5392
20101230,163300,1.5393,1.5394,1.5392,1.5392
20101230,163400,1.5391,1.5392,1.539,1.5392
20101230,163500,1.5391,1.5391,1.5391,1.5391
20101230,163600,1.5393,1.5393,1.5393,1.5393
20101230,163800,1.539,1.539,1.539,1.539
20101230,163900,1.5391,1.5391,1.5391,1.5391
20101230,164000,1.539,1.539,1.539,1.539
20101230,164200,1.5392,1.5392,1.5392,1.5392
20101230,164300,1.539,1.539,1.539,1.539
20101230,164400,1.5387,1.5387,1.5387,1.5387
20101230,164600,1.5386,1.5387,1.5384,1.5385
20101230,164700,1.5383,1.5383,1.5383,1.5383
20101230,164800,1.538,1.538,1.538,1.538
20101230,164900,1.5381,1.5381,1.5381,1.5381
20101230,165000,1.5383,1.5383,1.5383,1.5383
20101230,165100,1.5386,1.5386,1.5386,1.5386
20101230,165300,1.5385,1.5386,1.5384,1.5386
20101230,165400,1.5385,1.5385,1.5383,1.5383
20101230,165500,1.5382,1.5382,1.5381,1.5382
20101230,165600,1.5381,1.5386,1.5381,1.5382
20101230,165800,1.5394,1.5394,1.5394,1.5394
20101230,165900,1.5389,1.5389,1.5389,1.5389
20101230,170100,1.5388,1.5388,1.5381,1.5381
20101230,170200,1.5381,1.5381,1.5381,1.5381
20101230,170300,1.538,1.538,1.538,1.538
20101230,170400,1.5382,1.5382,1.5382,1.5382
20101230,170500,1.538,1.538,1.538,1.538
20101230,170600,1.5376,1.5376,1.5376,1.5376
20101230,170800,1.5377,1.5381,1.5376,1.5381
20101230,170900,1.5378,1.5378,1.5378,1.5378
20101230,171100,1.5375,1.5375,1.5375,1.5375
20101230,171200,1.5369,1.5369,1.5369,1.5369
20101230,171300,1.537,1.537,1.537,1.537
20101230,171500,1.537,1.537,1.537,1.537
20101230,171600,1.537,1.537,1.537,1.537
20101230,171700,1.5371,1.5371,1.5371,1.5371
20101230,171900,1.537,1.537,1.537,1.537
20101230,172000,1.537,1.537,1.537,1.537
20101230,172200,1.5369,1.5371,1.5369,1.537
20101230,172300,1.537,1.5372,1.537,1.5371
20101230,172400,1.5368,1.5368,1.5368,1.5368
20101230,172500,1.5366,1.5366,1.5366,1.5366
20101230,172600,1.5367,1.5367,1.5366,1.5367
20101230,172800,1.5367,1.5369,1.5367,1.5368
20101230,172900,1.5369,1.5374,1.5369,1.5374
20101230,173000,1.5374,1.5374,1.5374,1.5374
20101230,173100,1.5373,1.5373,1.5371,1.5371
20101230,173200,1.537,1.537,1.537,1.537
20101230,173400,1.5369,1.5369,1.5369,1.5369
20101230,173500,1.5371,1.5371,1.5371,1.5371
20101230,173700,1.5369,1.5369,1.5369,1.5369
20101230,173900,1.5369,1.5371,1.5369,1.5371
20101230,174000,1.5371,1.5371,1.5369,1.5369
20101230,174100,1.537,1.537,1.5369,1.5369
20101230,174200,1.5369,1.537,1.5367,1.5368
20101230,174300,1.5368,1.5368,1.5368,1.5368
20101230,174500,1.5368,1.5368,1.5368,1.5368
20101230,174600,1.5369,1.5369,1.5369,1.5369
20101230,174700,1.5372,1.5372,1.5372,1.5372
20101230,174900,1.5372,1.5373,1.5372,1.5373
20101230,175000,1.5372,1.5373,1.5372,1.5373
20101230,175100,1.5374,1.5374,1.5374,1.5374
20101230,175200,1.5374,1.5374,1.5374,1.5374
20101230,175300,1.5376,1.5376,1.5376,1.5376
20101230,175400,1.538,1.538,1.538,1.538
20101230,175500,1.5381,1.5381,1.5381,1.5381
20101230,175600,1.5385,1.5385,1.5385,1.5385
20101230,175800,1.5387,1.5387,1.5387,1.5387
20101230,180000,1.5387,1.5391,1.5385,1.5391
20101230,180100,1.5392,1.5392,1.5385,1.5385
20101230,180200,1.5386,1.5386,1.5385,1.5386
20101230,180300,1.5386,1.5386,1.5385,1.5385
20101230,180400,1.5385,1.5385,1.5384,1.5384
20101230,180500,1.5384,1.5385,1.5384,1.5385
20101230,180600,1.5384,1.5385,1.5384,1.5384
20101230,180700,1.5383,1.5385,1.5383,1.5385
20101230,180800,1.5384,1.5385,1.5384,1.5385
20101230,180900,1.5385,1.5385,1.5383,1.5383
20101230,181000,1.5384,1.5386,1.5384,1.5386
20101230,181100,1.5386,1.5388,1.5385,1.5386
20101230,181200,1.5385,1.5388,1.5385,1.5387
20101230,181300,1.5388,1.539,1.5387,1.539
20101230,181400,1.5391,1.5391,1.539,1.539
20101230,181500,1.539,1.539,1.5389,1.5389
20101230,181600,1.539,1.539,1.5389,1.5389
20101230,181700,1.539,1.539,1.539,1.539
20101230,181800,1.539,1.5393,1.539,1.5393
20101230,181900,1.5394,1.5398,1.5394,1.5398
20101230,182000,1.5399,1.5401,1.5399,1.54
20101230,182100,1.5401,1.5402,1.5398,1.5398
20101230,182200,1.5397,1.54,1.5397,1.5399
20101230,182300,1.54,1.5401,1.54,1.5401
20101230,182400,1.54,1.5402,1.54,1.5402
20101230,182500,1.5402,1.5407,1.5401,1.5407
20101230,182600,1.5408,1.5409,1.5408,1.5408
20101230,182700,1.5407,1.5413,1.5407,1.5412
20101230,182800,1.5411,1.5411,1.5407,1.5407
20101230,182900,1.5406,1.5406,1.5403,1.5403
20101230,183000,1.5402,1.5402,1.54,1.5401
20101230,183100,1.5402,1.5406,1.5402,1.5406
20101230,183200,1.5405,1.5407,1.5404,1.5407
20101230,183300,1.5407,1.5407,1.5405,1.5405
20101230,183400,1.5405,1.5406,1.5405,1.5406
20101230,183500,1.5407,1.541,1.5407,1.5407
20101230,183600,1.5407,1.5408,1.5406,1.5407
20101230,183700,1.5406,1.5408,1.5406,1.5407
20101230,183800,1.5407,1.5408,1.5406,1.5408
20101230,183900,1.5407,1.5407,1.5407,1.5407
20101230,184000,1.5407,1.5411,1.5407,1.5411
20101230,184100,1.5411,1.5413,1.5411,1.5412
20101230,184200,1.5411,1.5411,1.5408,1.5408
20101230,184300,1.5408,1.5408,1.5407,1.5407
20101230,184400,1.5407,1.541,1.5407,1.541
20101230,184500,1.541,1.5411,1.541,1.5411
20101230,184600,1.5411,1.5412,1.5411,1.5412
20101230,184700,1.5412,1.5412,1.541,1.541
20101230,184800,1.541,1.5411,1.541,1.5411
20101230,184900,1.5411,1.5411,1.541,1.5411
20101230,185000,1.5411,1.5412,1.5411,1.5412
20101230,185100,1.5411,1.5411,1.5411,1.5411
20101230,185200,1.541,1.5412,1.541,1.5412
20101230,185300,1.5412,1.5414,1.5412,1.5412
20101230,185400,1.5414,1.5414,1.5412,1.5412
20101230,185500,1.5413,1.5414,1.5413,1.5414
20101230,185600,1.5414,1.5416,1.5414,1.5415
20101230,185700,1.5416,1.5417,1.5415,1.5417
20101230,185800,1.5416,1.5418,1.5416,1.5418
20101230,185900,1.5419,1.5419,1.5419,1.5419
20101230,190000,1.5419,1.5419,1.5417,1.5418
20101230,190100,1.5417,1.5418,1.5416,1.5418
20101230,190200,1.5418,1.5418,1.5417,1.5417
20101230,190300,1.5417,1.5418,1.5417,1.5417
20101230,190400,1.5418,1.5421,1.5418,1.542
20101230,190500,1.542,1.542,1.5418,1.5418
20101230,190600,1.5418,1.5421,1.5417,1.5421
20101230,190700,1.5422,1.5423,1.5422,1.5422
20101230,190800,1.5422,1.5422,1.542,1.542
20101230,190900,1.542,1.542,1.5418,1.542
20101230,191000,1.5419,1.542,1.5418,1.5418
20101230,191100,1.5417,1.5419,1.5417,1.5419
20101230,191200,1.5419,1.5421,1.5419,1.5421
20101230,191300,1.5422,1.5422,1.5421,1.5421
20101230,191400,1.5421,1.5421,1.5419,1.5419
20101230,191500,1.5419,1.5425,1.5419,1.5425
20101230,191600,1.5426,1.5426,1.5425,1.5425
20101230,191700,1.5425,1.5428,1.5425,1.5428
20101230,191800,1.5429,1.5429,1.5428,1.5428
20101230,191900,1.5428,1.5428,1.5427,1.5428
20101230,192000,1.5428,1.5428,1.5425,1.5425
20101230,192100,1.5425,1.5425,1.5424,1.5424
20101230,192200,1.5424,1.5426,1.5424,1.5425
20101230,192300,1.5426,1.5428,1.5425,1.5425
20101230,192400,1.5425,1.5425,1.5423,1.5423
20101230,192500,1.5424,1.5424,1.542,1.5421
20101230,192600,1.5421,1.5422,1.5421,1.5421
20101230,192700,1.5421,1.5422,1.5421,1.5422
20101230,192800,1.5422,1.5422,1.5421,1.5422
20101230,192900,1.5421,1.5422,1.5421,1.5421
20101230,193000,1.5421,1.5421,1.542,1.542
20101230,193100,1.542,1.542,1.5419,1.542
20101230,193200,1.542,1.5422,1.5419,1.5422
20101230,193300,1.5422,1.5422,1.5422,1.5422
20101230,193400,1.5421,1.5421,1.5419,1.5419
20101230,193500,1.5419,1.542,1.5418,1.5419
20101230,193600,1.5418,1.5419,1.5418,1.5419
20101230,193700,1.5418,1.5419,1.5418,1.5418
20101230,193800,1.5419,1.542,1.5419,1.542
20101230,193900,1.5419,1.5421,1.5419,1.542
20101230,194000,1.5419,1.5423,1.5419,1.5423
20101230,194100,1.5422,1.5422,1.542,1.542
20101230,194200,1.5419,1.5422,1.5419,1.5422
20101230,194300,1.5423,1.5424,1.5422,1.5422
20101230,194400,1.5422,1.5422,1.542,1.5421
20101230,194500,1.542,1.5422,1.542,1.5422
20101230,194600,1.5423,1.5423,1.5423,1.5423
20101230,194700,1.5422,1.5422,1.5421,1.5421
20101230,194800,1.5421,1.5422,1.5421,1.5422
20101230,194900,1.5421,1.5422,1.542,1.5422
20101230,195000,1.5421,1.5421,1.5418,1.5418
20101230,195100,1.5418,1.5419,1.5417,1.5418
20101230,195200,1.5417,1.5418,1.5417,1.5418
20101230,195300,1.5419,1.5419,1.5417,1.5418
20101230,195400,1.5417,1.5418,1.5417,1.5418
20101230,195500,1.5418,1.5418,1.5414,1.5414
20101230,195600,1.5415,1.5415,1.5415,1.5415
20101230,195700,1.5415,1.5416,1.5415,1.5416
20101230,195800,1.5415,1.5416,1.5414,1.5414
20101230,195900,1.5414,1.5414,1.5411,1.5411
20101230,200000,1.5412,1.5413,1.5412,1.5413
20101230,200100,1.5413,1.5414,1.5412,1.5412
20101230,200200,1.5413,1.5413,1.541,1.541
20101230,200300,1.5411,1.5411,1.5408,1.5408
20101230,200400,1.5408,1.5409,1.5408,1.5409
20101230,200500,1.5409,1.541,1.5408,1.5409
20101230,200600,1.5409,1.541,1.5409,1.5409
20101230,200700,1.541,1.5411,1.5409,1.541
20101230,200800,1.541,1.541,1.541,1.541
20101230,200900,1.5409,1.541,1.5409,1.5409
20101230,201000,1.5409,1.541,1.5408,1.541
20101230,201100,1.5411,1.5411,1.5409,1.5411
20101230,201200,1.5411,1.5412,1.5411,1.5412
20101230,201300,1.5413,1.5414,1.5413,1.5414
20101230,201400,1.5414,1.5414,1.5413,1.5413
20101230,201500,1.5414,1.5415,1.5414,1.5415
20101230,201600,1.5415,1.5415,1.5414,1.5414
20101230,201700,1.5414,1.5415,1.5414,1.5414
20101230,201800,1.5413,1.5413,1.5412,1.5413
20101230,201900,1.5413,1.5415,1.5413,1.5415
20101230,202000,1.5415,1.5416,1.5415,1.5416
20101230,202100,1.5416,1.5417,1.5416,1.5417
20101230,202200,1.5417,1.5419,1.5417,1.5419
20101230,202300,1.542,1.542,1.5418,1.5418
20101230,202400,1.5418,1.5419,1.5418,1.5419
20101230,202500,1.5418,1.5419,1.5418,1.5419
20101230,202600,1.5418,1.5419,1.5417,1.5419
20101230,202700,1.5418,1.5419,1.5418,1.5419
20101230,202800,1.5419,1.5419,1.5417,1.5417
20101230,202900,1.5417,1.5417,1.5416,1.5416
20101230,203000,1.5416,1.5416,1.5415,1.5415
20101230,203100,1.5416,1.5419,1.5416,1.5419
20101230,203200,1.5418,1.5421,1.5417,1.5421
20101230,203300,1.5421,1.5421,1.542,1.5421
20101230,203400,1.5421,1.5421,1.5419,1.5421
20101230,203500,1.5421,1.5421,1.542,1.5421
20101230,203600,1.5421,1.5421,1.5419,1.5419
20101230,203700,1.5418,1.5419,1.5416,1.5416
20101230,203800,1.5416,1.5416,1.5414,1.5416
20101230,203900,1.5416,1.5416,1.5416,1.5416
20101230,204000,1.5416,1.5417,1.5416,1.5417
20101230,204100,1.5416,1.5416,1.5415,1.5416
20101230,204200,1.5415,1.5416,1.5415,1.5415
20101230,204300,1.5414,1.5414,1.5414,1.5414
20101230,204400,1.5414,1.5414,1.5412,1.5412
20101230,204500,1.5412,1.5412,1.5412,1.5412
20101230,204600,1.5412,1.5412,1.5411,1.5411
20101230,204700,1.5411,1.5412,1.5411,1.5411
20101230,204800,1.5411,1.5413,1.5411,1.5413
20101230,204900,1.5414,1.5414,1.5412,1.5414
20101230,205000,1.5413,1.5413,1.5413,1.5413
20101230,205100,1.5413,1.5413,1.5413,1.5413
20101230,205200,1.5413,1.5414,1.5412,1.5414
20101230,205300,1.5414,1.5415,1.5414,1.5415
20101230,205400,1.5414,1.5416,1.5413,1.5416
20101230,205500,1.5416,1.5417,1.5415,1.5417
20101230,205600,1.5417,1.5419,1.5417,1.5419
20101230,205700,1.542,1.5421,1.542,1.5421
20101230,205800,1.5421,1.5421,1.5419,1.5419
20101230,205900,1.5421,1.5421,1.5418,1.542
20101230,210000,1.5419,1.5421,1.5419,1.542
20101230,210100,1.5419,1.5419,1.5418,1.5419
20101230,210200,1.542,1.5421,1.542,1.542
20101230,210300,1.5421,1.5422,1.5421,1.5422
20101230,210400,1.542,1.5423,1.542,1.5423
20101230,210500,1.5423,1.5424,1.5423,1.5424
20101230,210600,1.5423,1.5424,1.5422,1.5422
20101230,210700,1.5421,1.5424,1.5421,1.5423
20101230,210800,1.5423,1.5423,1.5421,1.5421
20101230,210900,1.5422,1.5422,1.542,1.542
20101230,211000,1.5421,1.5421,1.542,1.5421
20101230,211100,1.5419,1.542,1.5418,1.5418
20101230,211200,1.5419,1.5421,1.5419,1.5419
20101230,211300,1.5418,1.5419,1.5418,1.5419
20101230,211400,1.5419,1.542,1.5419,1.542
20101230,211500,1.542,1.542,1.542,1.542
20101230,211600,1.542,1.542,1.5418,1.542
20101230,211700,1.5421,1.5421,1.5417,1.542
20101230,211800,1.5421,1.5421,1.5418,1.5418
20101230,211900,1.5417,1.5417,1.5417,1.5417
20101230,212000,1.5416,1.5418,1.5416,1.5418
20101230,212100,1.5418,1.5419,1.5418,1.5418
20101230,212200,1.5418,1.5419,1.5417,1.5418
20101230,212300,1.5419,1.542,1.5418,1.5418
20101230,212400,1.5419,1.5421,1.5418,1.5421
20101230,212500,1.5421,1.5421,1.542,1.542
20101230,212600,1.5419,1.542,1.5418,1.542
20101230,212700,1.542,1.5423,1.542,1.5421
20101230,212800,1.5421,1.5423,1.542,1.5423
20101230,212900,1.5424,1.5424,1.5422,1.5424
20101230,213000,1.5423,1.5423,1.5422,1.5423
20101230,213100,1.5423,1.5423,1.5423,1.5423
20101230,213200,1.5422,1.5423,1.542,1.5423
20101230,213300,1.5423,1.5426,1.5422,1.5424
20101230,213400,1.5425,1.5425,1.5423,1.5425
20101230,213500,1.5426,1.5426,1.5423,1.5426
20101230,213600,1.5425,1.5427,1.5423,1.5423
20101230,213700,1.5424,1.5424,1.5424,1.5424
20101230,213800,1.5424,1.5424,1.5422,1.5423
20101230,213900,1.5424,1.5424,1.5422,1.5423
20101230,214000,1.5423,1.5424,1.5423,1.5423
20101230,214100,1.5422,1.5422,1.5421,1.5421
20101230,214200,1.5422,1.5423,1.5422,1.5423
20101230,214300,1.5423,1.5424,1.5423,1.5423
20101230,214400,1.5423,1.5423,1.5423,1.5423
20101230,214500,1.5423,1.5423,1.5423,1.5423
20101230,214600,1.5424,1.5424,1.5423,1.5423
20101230,214700,1.5423,1.5424,1.5423,1.5423
20101230,214800,1.5424,1.5424,1.5423,1.5424
20101230,214900,1.5423,1.5423,1.5423,1.5423
20101230,215000,1.5423,1.5423,1.5422,1.5423
20101230,215100,1.5423,1.5424,1.5422,1.5424
20101230,215200,1.5424,1.5424,1.5424,1.5424
20101230,215300,1.5424,1.5424,1.5424,1.5424
20101230,215400,1.5424,1.5424,1.5424,1.5424
20101230,215500,1.5423,1.5424,1.5423,1.5423
20101230,215600,1.5423,1.5423,1.5423,1.5423
20101230,215700,1.5424,1.5424,1.5423,1.5424
20101230,215800,1.5424,1.5424,1.5424,1.5424
20101230,215900,1.5424,1.5424,1.5423,1.5423
20101230,220000,1.5424,1.5425,1.5424,1.5424
20101230,220100,1.5425,1.5427,1.5424,1.5427
20101230,220200,1.5426,1.5426,1.5424,1.5425
20101230,220300,1.5425,1.5425,1.5425,1.5425
20101230,220400,1.5426,1.5426,1.5425,1.5425
20101230,220500,1.5425,1.5425,1.5423,1.5423
20101230,220600,1.5423,1.5424,1.5423,1.5424
20101230,220700,1.5425,1.5426,1.5423,1.5423
20101230,220800,1.5424,1.5425,1.5424,1.5425
20101230,220900,1.5425,1.5427,1.5425,1.5427
20101230,221000,1.5427,1.5427,1.5425,1.5425
20101230,221100,1.5426,1.5426,1.5425,1.5425
20101230,221200,1.5425,1.5426,1.5425,1.5426
20101230,221300,1.5425,1.5425,1.5424,1.5424
20101230,221400,1.5424,1.5425,1.5424,1.5424
20101230,221500,1.5425,1.5425,1.5425,1.5425
20101230,221600,1.5426,1.5426,1.5426,1.5426
20101230,221700,1.5426,1.5426,1.5425,1.5425
20101230,221800,1.5426,1.5426,1.5425,1.5425
20101230,221900,1.5425,1.5426,1.5425,1.5426
20101230,222000,1.5425,1.5425,1.5425,1.5425
20101230,222100,1.5425,1.5426,1.5424,1.5424
20101230,222200,1.5424,1.5424,1.5424,1.5424
20101230,222300,1.5423,1.5426,1.5423,1.5426
20101230,222400,1.5426,1.5426,1.5423,1.5426
20101230,222500,1.5425,1.5425,1.5424,1.5425
20101230,222600,1.5425,1.5425,1.5423,1.5425
20101230,222700,1.5425,1.5427,1.5425,1.5426
20101230,222800,1.5426,1.5426,1.5425,1.5425
20101230,222900,1.5425,1.5426,1.5425,1.5426
20101230,223000,1.5425,1.5426,1.5425,1.5426
20101230,223100,1.5426,1.5426,1.5426,1.5426
20101230,223200,1.5425,1.5425,1.5425,1.5425
20101230,223300,1.5424,1.5425,1.5424,1.5424
20101230,223400,1.5424,1.5424,1.5423,1.5423
20101230,223500,1.5423,1.5424,1.5423,1.5424
20101230,223600,1.5424,1.5424,1.5423,1.5423
20101230,223700,1.5423,1.5425,1.5423,1.5425
20101230,223800,1.5425,1.5426,1.5425,1.5426
20101230,223900,1.5425,1.5425,1.5424,1.5424
20101230,224000,1.5424,1.5424,1.5423,1.5423
20101230,224100,1.5423,1.5424,1.5423,1.5424
20101230,224200,1.5424,1.5425,1.5424,1.5425
20101230,224300,1.5425,1.5425,1.5425,1.5425
20101230,224400,1.5425,1.5426,1.5425,1.5426
20101230,224500,1.5426,1.5426,1.5426,1.5426
20101230,224600,1.5426,1.5426,1.5426,1.5426
20101230,224700,1.5426,1.5427,1.5426,1.5427
20101230,224800,1.5429,1.5429,1.5429,1.5429
20101230,224900,1.5427,1.5427,1.5427,1.5427
20101230,225100,1.5427,1.5427,1.5427,1.5427
20101230,225200,1.5427,1.5427,1.5427,1.5427
20101230,225400,1.5427,1.5427,1.5425,1.5426
20101230,225500,1.5426,1.5426,1.5426,1.5426
20101230,225700,1.5426,1.5426,1.5426,1.5426
20101230,225800,1.5426,1.5426,1.5426,1.5426
20101230,225900,1.5428,1.5428,1.5428,1.5428
20101230,230100,1.5431,1.5431,1.5431,1.5431
20101230,230200,1.5432,1.5432,1.5432,1.5432
20101230,230300,1.5432,1.5432,1.5432,1.5432
20101230,230400,1.5432,1.5432,1.5432,1.5432
20101230,230500,1.543,1.543,1.543,1.543
20101230,230700,1.5429,1.5429,1.5429,1.5429
20101230,230900,1.543,1.5431,1.543,1.5431
20101230,231000,1.5433,1.5433,1.5433,1.5433
20101230,231200,1.5431,1.5431,1.5431,1.5431
20101230,231400,1.5428,1.5428,1.5428,1.5428
20101230,231500,1.5427,1.5427,1.5427,1.5427
20101230,231600,1.5423,1.5423,1.5423,1.5423
20101230,231700,1.5426,1.5426,1.5426,1.5426
20101230,231900,1.5427,1.5427,1.5427,1.5427
20101230,232100,1.5427,1.5427,1.5425,1.5425
20101230,232200,1.5426,1.5426,1.5426,1.5426
20101230,232300,1.5425,1.5425,1.5425,1.5425
20101230,232400,1.5424,1.5424,1.5424,1.5424
20101230,232500,1.5427,1.5427,1.5427,1.5427
20101230,232700,1.5425,1.5425,1.5425,1.5425
20101230,232900,1.5426,1.5426,1.5426,1.5426
20101230,233000,1.5426,1.5426,1.5426,1.5426
20101230,233200,1.5428,1.5428,1.5428,1.5428
20101230,233300,1.5427,1.5427,1.5427,1.5427
20101230,233400,1.5425,1.5425,1.5425,1.5425
20101230,233600,1.5428,1.5428,1.5428,1.5428
20101230,233800,1.5427,1.5428,1.5426,1.5428
20101230,233900,1.5432,1.5432,1.543,1.543
20101230,234000,1.5431,1.5432,1.5431,1.5431
20101230,234100,1.5432,1.5432,1.5429,1.543
20101230,234200,1.543,1.5431,1.543,1.543
20101230,234300,1.543,1.543,1.543,1.543
20101230,234400,1.543,1.543,1.5428,1.5429
20101230,234500,1.5431,1.5431,1.5431,1.5431
20101230,234600,1.5432,1.5432,1.543,1.543
20101230,234700,1.5431,1.5431,1.543,1.543
20101230,234800,1.543,1.5432,1.5428,1.543
20101230,235000,1.5432,1.5432,1.543,1.543
20101230,235100,1.543,1.543,1.543,1.543
20101230,235200,1.543,1.543,1.5428,1.5428
20101230,235300,1.5428,1.543,1.5428,1.543
20101230,235400,1.5432,1.5432,1.5432,1.5432
20101230,235600,1.5433,1.5433,1.5433,1.5433
20101230,235700,1.5433,1.5435,1.5433,1.5433
20101230,235900,1.5433,1.5435,1.5433,1.5435
20101231,0,1.5433,1.5434,1.5433,1.5433
20101231,100,1.5433,1.5433,1.5433,1.5433
20101231,200,1.5436,1.5436,1.5432,1.5432
20101231,300,1.5432,1.5432,1.5431,1.5431
20101231,400,1.5431,1.5432,1.5431,1.5432
20101231,500,1.5431,1.5433,1.5431,1.5433
20101231,600,1.5432,1.5433,1.5431,1.5433
20101231,700,1.5434,1.5434,1.5432,1.5433
20101231,800,1.5431,1.5435,1.5431,1.5433
20101231,900,1.5433,1.5433,1.5431,1.5431
20101231,1000,1.5431,1.5433,1.5431,1.5433
20101231,1100,1.5432,1.5434,1.5432,1.5434
20101231,1200,1.5433,1.5434,1.5432,1.5432
20101231,1300,1.5432,1.5432,1.5431,1.5431
20101231,1400,1.5432,1.5434,1.5432,1.5433
20101231,1500,1.5434,1.5434,1.5434,1.5434
20101231,1600,1.5434,1.5434,1.5433,1.5434
20101231,1700,1.5434,1.5435,1.5432,1.5432
20101231,1800,1.5432,1.5434,1.5432,1.5434
20101231,1900,1.5435,1.5435,1.5432,1.5432
20101231,2000,1.5432,1.5434,1.5432,1.5432
20101231,2100,1.5432,1.5434,1.5432,1.5434
20101231,2200,1.5434,1.5434,1.5432,1.5432
20101231,2300,1.5433,1.5433,1.543,1.543
20101231,2400,1.5431,1.5432,1.543,1.5431
20101231,2500,1.543,1.5432,1.543,1.5432
20101231,2600,1.5432,1.5433,1.5432,1.5433
20101231,2700,1.5432,1.5433,1.5431,1.5431
20101231,2800,1.5432,1.5432,1.5432,1.5432
20101231,2900,1.5432,1.5432,1.5432,1.5432
20101231,3000,1.5432,1.5433,1.5432,1.5433
20101231,3100,1.5434,1.5434,1.5433,1.5433
20101231,3200,1.5434,1.5434,1.5431,1.5432
20101231,3300,1.5432,1.5432,1.5431,1.5432
20101231,3400,1.5432,1.5433,1.5432,1.5432
20101231,3500,1.5432,1.5434,1.5432,1.5433
20101231,3600,1.5433,1.5435,1.5433,1.5435
20101231,3700,1.5435,1.5435,1.5433,1.5433
20101231,3800,1.5434,1.5434,1.5433,1.5433
20101231,3900,1.5433,1.5434,1.5433,1.5434
20101231,4000,1.5433,1.5434,1.5433,1.5434
20101231,4100,1.5434,1.5435,1.543,1.5431
20101231,4200,1.5431,1.5433,1.5431,1.5432
20101231,4300,1.5431,1.5431,1.543,1.543
20101231,4400,1.5431,1.5431,1.543,1.5431
20101231,4500,1.5431,1.5433,1.5431,1.5433
20101231,4600,1.5432,1.5432,1.5431,1.5431
20101231,4700,1.5431,1.5433,1.5431,1.5432
20101231,4800,1.5432,1.5432,1.5427,1.5427
20101231,4900,1.5426,1.5427,1.5426,1.5427
20101231,5000,1.5427,1.5428,1.5426,1.5426
20101231,5100,1.5426,1.5426,1.5426,1.5426
20101231,5200,1.5425,1.5425,1.5424,1.5425
20101231,5300,1.5424,1.5424,1.5423,1.5423
20101231,5400,1.5424,1.5425,1.5424,1.5425
20101231,5500,1.5426,1.5432,1.5426,1.543
20101231,5600,1.5431,1.5433,1.5431,1.5433
20101231,5700,1.5433,1.5434,1.5433,1.5434
20101231,5800,1.5435,1.5435,1.5435,1.5435
20101231,5900,1.5436,1.5436,1.5435,1.5435
20101231,10000,1.5435,1.5435,1.5431,1.5433
20101231,10100,1.5432,1.5435,1.5432,1.5435
20101231,10200,1.5436,1.5436,1.5434,1.5434
20101231,10300,1.5434,1.5436,1.5434,1.5436
20101231,10400,1.5436,1.5437,1.5436,1.5436
20101231,10500,1.5436,1.5437,1.5436,1.5437
20101231,10600,1.5438,1.544,1.5437,1.5439
20101231,10700,1.5439,1.544,1.5438,1.544
20101231,10800,1.544,1.5441,1.5439,1.5441
20101231,10900,1.5441,1.5441,1.544,1.5441
20101231,11000,1.544,1.5441,1.5439,1.5441
20101231,11100,1.5441,1.5441,1.5441,1.5441
20101231,11200,1.544,1.5441,1.5439,1.544
20101231,11300,1.5441,1.5442,1.5441,1.5442
20101231,11400,1.5441,1.5441,1.544,1.544
20101231,11500,1.544,1.5441,1.544,1.5441
20101231,11600,1.5441,1.5445,1.5441,1.5444
20101231,11700,1.5444,1.5445,1.5444,1.5445
20101231,11800,1.5444,1.5444,1.5443,1.5443
20101231,11900,1.5443,1.5444,1.5443,1.5444
20101231,12000,1.5444,1.5444,1.5443,1.5444
20101231,12100,1.5443,1.5444,1.5442,1.5444
20101231,12200,1.5444,1.5444,1.5442,1.5443
20101231,12300,1.5443,1.5444,1.5443,1.5444
20101231,12400,1.5444,1.5444,1.5442,1.5442
20101231,12500,1.5442,1.5444,1.5442,1.5444
20101231,12600,1.5444,1.5444,1.5442,1.5444
20101231,12700,1.5444,1.5444,1.5443,1.5443
20101231,12800,1.5443,1.5443,1.5443,1.5443
20101231,12900,1.5443,1.5443,1.5443,1.5443
20101231,13000,1.5443,1.5444,1.5441,1.5441
20101231,13100,1.544,1.5441,1.5439,1.5441
20101231,13200,1.5441,1.5441,1.5441,1.5441
20101231,13300,1.5442,1.5442,1.544,1.544
20101231,13400,1.544,1.5442,1.5439,1.5442
20101231,13500,1.5442,1.5442,1.5441,1.5441
20101231,13600,1.5442,1.5443,1.5442,1.5442
20101231,13700,1.544,1.5441,1.544,1.544
20101231,13800,1.544,1.5442,1.544,1.5442
20101231,13900,1.5442,1.5442,1.5441,1.5442
20101231,14000,1.544,1.544,1.5438,1.544
20101231,14100,1.544,1.5443,1.544,1.5442
20101231,14200,1.5442,1.5442,1.544,1.5441
20101231,14300,1.544,1.5443,1.544,1.5441
20101231,14400,1.5441,1.5442,1.544,1.5442
20101231,14500,1.5441,1.5441,1.544,1.5441
20101231,14600,1.5441,1.5441,1.544,1.5441
20101231,14700,1.544,1.5441,1.5437,1.5437
20101231,14800,1.5438,1.5439,1.5438,1.5439
20101231,14900,1.544,1.544,1.5438,1.5438
20101231,15000,1.5438,1.5439,1.5435,1.5439
20101231,15100,1.5438,1.5439,1.5438,1.5439
20101231,15200,1.5439,1.5439,1.5435,1.5435
20101231,15300,1.5435,1.5438,1.5435,1.5438
20101231,15400,1.5439,1.544,1.5439,1.544
20101231,15500,1.5439,1.5441,1.5439,1.5441
20101231,15600,1.5441,1.5441,1.5441,1.5441
20101231,15700,1.5441,1.5441,1.5441,1.5441
20101231,15800,1.5441,1.5441,1.5441,1.5441
20101231,15900,1.5441,1.5442,1.544,1.5441
20101231,20000,1.544,1.5441,1.544,1.5441
20101231,20100,1.5441,1.5442,1.5441,1.5441
20101231,20200,1.5441,1.5442,1.544,1.5442
20101231,20300,1.5441,1.5441,1.544,1.5441
20101231,20400,1.5441,1.5441,1.5441,1.5441
20101231,20500,1.5441,1.5441,1.5439,1.544
20101231,20600,1.5441,1.5441,1.5439,1.5441
20101231,20700,1.5442,1.5443,1.5442,1.5443
20101231,20800,1.5444,1.5446,1.5444,1.5446
20101231,20900,1.5445,1.5446,1.5444,1.5445
20101231,21000,1.5446,1.5446,1.5445,1.5445
20101231,21100,1.5446,1.5453,1.5445,1.5453
20101231,21200,1.5453,1.5453,1.5453,1.5453
20101231,21300,1.5453,1.5454,1.5453,1.5453
20101231,21400,1.5452,1.5452,1.5451,1.5452
20101231,21500,1.5452,1.5452,1.545,1.5451
20101231,21600,1.5452,1.5452,1.5452,1.5452
20101231,21700,1.545,1.5454,1.545,1.5454
20101231,21800,1.5455,1.5459,1.5455,1.5459
20101231,21900,1.5458,1.5459,1.5457,1.5458
20101231,22000,1.5457,1.5459,1.5457,1.5459
20101231,22100,1.5458,1.5459,1.5456,1.5456
20101231,22200,1.5457,1.5458,1.5456,1.5456
20101231,22300,1.5455,1.5456,1.5454,1.5456
20101231,22400,1.5455,1.5456,1.5453,1.5455
20101231,22500,1.5456,1.5456,1.5452,1.5454
20101231,22600,1.5454,1.5454,1.5453,1.5453
20101231,22700,1.5452,1.5453,1.5452,1.5452
20101231,22800,1.5451,1.5452,1.5447,1.5448
20101231,22900,1.5447,1.5448,1.5446,1.5447
20101231,23000,1.5448,1.5448,1.5447,1.5447
20101231,23100,1.5446,1.5446,1.5445,1.5446
20101231,23200,1.5445,1.5445,1.5444,1.5445
20101231,23300,1.5443,1.5446,1.5443,1.5444
20101231,23400,1.5444,1.5445,1.5444,1.5445
20101231,23500,1.5444,1.5445,1.5442,1.5445
20101231,23600,1.5444,1.5445,1.5443,1.5443
20101231,23700,1.5442,1.5446,1.5442,1.5445
20101231,23800,1.5446,1.545,1.5446,1.5449
20101231,23900,1.545,1.545,1.5449,1.5449
20101231,24000,1.5449,1.545,1.5448,1.5449
20101231,24100,1.5447,1.5451,1.5447,1.5451
20101231,24200,1.545,1.5451,1.545,1.545
20101231,24300,1.5449,1.545,1.5448,1.5448
20101231,24400,1.5448,1.545,1.5448,1.545
20101231,24500,1.545,1.545,1.5449,1.5449
20101231,24600,1.5449,1.545,1.5449,1.545
20101231,24700,1.545,1.5451,1.545,1.545
20101231,24800,1.5449,1.5449,1.5445,1.5447
20101231,24900,1.5448,1.5448,1.5448,1.5448
20101231,25000,1.5448,1.5448,1.5446,1.5447
20101231,25100,1.5447,1.5448,1.5446,1.5448
20101231,25200,1.5447,1.5447,1.5444,1.5444
20101231,25300,1.5443,1.5444,1.5442,1.5442
20101231,25400,1.5442,1.5446,1.5441,1.5445
20101231,25500,1.5444,1.5444,1.5443,1.5443
20101231,25600,1.5442,1.5444,1.5442,1.5444
20101231,25700,1.5443,1.5444,1.5443,1.5444
20101231,25800,1.5445,1.5446,1.5445,1.5445
20101231,25900,1.5445,1.5445,1.5441,1.5441
20101231,30000,1.5441,1.5441,1.544,1.5441
20101231,30100,1.5441,1.5442,1.544,1.5441
20101231,30200,1.5442,1.5442,1.5441,1.5441
20101231,30300,1.5441,1.5444,1.544,1.5444
20101231,30400,1.5445,1.5445,1.5442,1.5442
20101231,30500,1.5442,1.5444,1.5442,1.5443
20101231,30600,1.5442,1.5443,1.5442,1.5442
20101231,30700,1.5441,1.5443,1.5441,1.5441
20101231,30800,1.5441,1.5444,1.5441,1.5444
20101231,30900,1.5445,1.5447,1.5445,1.5446
20101231,31000,1.5447,1.5447,1.5446,1.5447
20101231,31100,1.5447,1.5447,1.5447,1.5447
20101231,31200,1.5446,1.5446,1.5446,1.5446
20101231,31300,1.5446,1.5446,1.5446,1.5446
20101231,31400,1.5445,1.5449,1.5445,1.5449
20101231,31500,1.5448,1.5448,1.5447,1.5448
20101231,31600,1.5447,1.545,1.5447,1.545
20101231,31700,1.5449,1.5449,1.5448,1.5448
20101231,31800,1.5448,1.5448,1.5447,1.5448
20101231,31900,1.5447,1.5448,1.5447,1.5448
20101231,32000,1.5448,1.5448,1.5447,1.5447
20101231,32100,1.5447,1.5447,1.5446,1.5446
20101231,32200,1.5447,1.5447,1.5444,1.5444
20101231,32300,1.5445,1.5445,1.5444,1.5445
20101231,32400,1.5445,1.5445,1.5444,1.5444
20101231,32500,1.5443,1.5444,1.5441,1.5442
20101231,32600,1.5441,1.5442,1.5441,1.5441
20101231,32700,1.5442,1.5442,1.544,1.5441
20101231,32800,1.544,1.5441,1.544,1.5441
20101231,32900,1.5441,1.5441,1.5438,1.5439
20101231,33000,1.5438,1.5438,1.5432,1.5432
20101231,33100,1.5431,1.5433,1.5431,1.5433
20101231,33200,1.5434,1.5436,1.5432,1.5434
20101231,33300,1.5434,1.5434,1.5434,1.5434
20101231,33400,1.5433,1.5435,1.5433,1.5435
20101231,33500,1.5435,1.5436,1.5434,1.5435
20101231,33600,1.5434,1.5439,1.5434,1.5438
20101231,33700,1.5437,1.5437,1.5434,1.5435
20101231,33800,1.5433,1.5434,1.5433,1.5434
20101231,33900,1.5435,1.5435,1.5434,1.5435
20101231,34000,1.5435,1.5438,1.5435,1.5438
20101231,34100,1.5439,1.5439,1.5437,1.5437
20101231,34200,1.5438,1.5441,1.5438,1.5441
20101231,34300,1.5441,1.5443,1.544,1.544
20101231,34400,1.5439,1.544,1.5436,1.5437
20101231,34500,1.5438,1.5439,1.5438,1.5439
20101231,34600,1.544,1.544,1.5438,1.5439
20101231,34700,1.544,1.544,1.5439,1.5439
20101231,34800,1.5439,1.5439,1.5438,1.5439
20101231,34900,1.544,1.5443,1.544,1.5443
20101231,35000,1.5442,1.5442,1.5441,1.5441
20101231,35100,1.5442,1.5442,1.5441,1.5441
20101231,35200,1.5442,1.5442,1.5442,1.5442
20101231,35300,1.5442,1.5442,1.5439,1.5441
20101231,35400,1.5441,1.5441,1.5441,1.5441
20101231,35500,1.5442,1.5442,1.544,1.5441
20101231,35600,1.5441,1.5441,1.5439,1.5439
20101231,35700,1.5441,1.5441,1.5441,1.5441
20101231,35800,1.5441,1.5441,1.5441,1.5441
20101231,35900,1.5441,1.5441,1.5441,1.5441
20101231,40000,1.5441,1.5441,1.544,1.544
20101231,40100,1.5439,1.5443,1.5439,1.5443
20101231,40200,1.5442,1.5442,1.5438,1.5439
20101231,40300,1.544,1.5442,1.5439,1.5442
20101231,40400,1.5442,1.5442,1.5441,1.5441
20101231,40500,1.5442,1.5442,1.5438,1.5438
20101231,40600,1.5438,1.544,1.5438,1.544
20101231,40700,1.5441,1.5441,1.5435,1.5435
20101231,40800,1.5434,1.5435,1.5433,1.5435
20101231,40900,1.5436,1.5437,1.5435,1.5435
20101231,41000,1.5435,1.5435,1.5435,1.5435
20101231,41100,1.5436,1.5436,1.5435,1.5436
20101231,41200,1.5436,1.5436,1.5436,1.5436
20101231,41300,1.5437,1.5439,1.5437,1.5439
20101231,41400,1.5438,1.5438,1.5437,1.5438
20101231,41500,1.5438,1.5438,1.5436,1.5436
20101231,41600,1.5436,1.5436,1.5435,1.5435
20101231,41700,1.5436,1.5438,1.5436,1.5438
20101231,41800,1.5437,1.5438,1.5437,1.5437
20101231,41900,1.5438,1.5438,1.5438,1.5438
20101231,42000,1.5438,1.5438,1.5436,1.5436
20101231,42100,1.5437,1.5439,1.5437,1.5439
20101231,42200,1.5439,1.5439,1.5437,1.5439
20101231,42300,1.5438,1.5439,1.5438,1.5439
20101231,42400,1.5439,1.544,1.5438,1.5438
20101231,42500,1.5438,1.5438,1.5438,1.5438
20101231,42600,1.5438,1.5438,1.5437,1.5438
20101231,42700,1.5437,1.5438,1.5435,1.5435
20101231,42800,1.5436,1.5438,1.5436,1.5438
20101231,42900,1.5438,1.5439,1.5437,1.5439
20101231,43000,1.5438,1.5438,1.5438,1.5438
20101231,43100,1.5438,1.5439,1.5437,1.5438
20101231,43200,1.5438,1.5438,1.5436,1.5436
20101231,43300,1.5437,1.5437,1.5435,1.5437
20101231,43400,1.5436,1.5437,1.5436,1.5437
20101231,43500,1.5437,1.5437,1.5437,1.5437
20101231,43600,1.5437,1.5437,1.5437,1.5437
20101231,43700,1.5437,1.5437,1.5437,1.5437
20101231,43800,1.5437,1.5437,1.5436,1.5437
20101231,43900,1.5436,1.5437,1.5436,1.5437
20101231,44000,1.5436,1.5436,1.5436,1.5436
20101231,44100,1.5436,1.5437,1.5436,1.5437
20101231,44200,1.5437,1.5437,1.5436,1.5436
20101231,44300,1.5436,1.5438,1.5436,1.5437
20101231,44400,1.5437,1.5437,1.5435,1.5436
20101231,44500,1.5435,1.5435,1.5435,1.5435
20101231,44600,1.5434,1.5435,1.5432,1.5435
20101231,44700,1.5436,1.5439,1.5436,1.5437
20101231,44800,1.5436,1.5436,1.5436,1.5436
20101231,44900,1.5436,1.5438,1.5436,1.5438
20101231,45000,1.5437,1.5437,1.5437,1.5437
20101231,45100,1.5437,1.5438,1.5437,1.5438
20101231,45200,1.5437,1.5438,1.5437,1.5437
20101231,45300,1.5438,1.5439,1.5438,1.5439
20101231,45400,1.5439,1.5439,1.5437,1.5438
20101231,45500,1.5438,1.5439,1.5437,1.5439
20101231,45600,1.5439,1.544,1.5439,1.544
20101231,45700,1.544,1.544,1.5438,1.5438
20101231,45800,1.5439,1.5439,1.5437,1.5437
20101231,45900,1.5438,1.5438,1.5436,1.5436
20101231,50000,1.5437,1.5438,1.5432,1.5432
20101231,50100,1.5433,1.5435,1.5432,1.5434
20101231,50200,1.5434,1.5435,1.5434,1.5435
20101231,50300,1.5434,1.5434,1.5433,1.5434
20101231,50400,1.5434,1.5434,1.5433,1.5433
20101231,50500,1.5433,1.5433,1.5432,1.5432
20101231,50600,1.5433,1.5434,1.5432,1.5434
20101231,50700,1.5433,1.5434,1.5433,1.5434
20101231,50800,1.5433,1.5434,1.5433,1.5434
20101231,50900,1.5433,1.5433,1.5432,1.5433
20101231,51000,1.5433,1.5433,1.5433,1.5433
20101231,51100,1.5433,1.5434,1.5433,1.5433
20101231,51200,1.5432,1.5432,1.543,1.543
20101231,51300,1.5431,1.5432,1.5431,1.5432
20101231,51400,1.5431,1.5432,1.543,1.5432
20101231,51500,1.5433,1.5433,1.5431,1.5431
20101231,51600,1.5432,1.5437,1.5432,1.5436
20101231,51700,1.5434,1.5434,1.5433,1.5433
20101231,51800,1.5434,1.5435,1.5433,1.5433
20101231,51900,1.5434,1.5434,1.5434,1.5434
20101231,52000,1.5434,1.5434,1.5433,1.5433
20101231,52100,1.5431,1.5435,1.5431,1.5435
20101231,52200,1.5434,1.5436,1.5434,1.5435
20101231,52300,1.5434,1.5434,1.5432,1.5432
20101231,52400,1.5434,1.5435,1.5434,1.5435
20101231,52500,1.5434,1.5436,1.5434,1.5436
20101231,52600,1.5436,1.5436,1.5436,1.5436
20101231,52700,1.5437,1.5437,1.5436,1.5436
20101231,52800,1.5437,1.5439,1.5437,1.5437
20101231,52900,1.5437,1.5438,1.5437,1.5437
20101231,53000,1.5438,1.544,1.5438,1.5439
20101231,53100,1.5439,1.544,1.5437,1.544
20101231,53200,1.5439,1.5443,1.5439,1.5443
20101231,53300,1.5443,1.5443,1.5441,1.5441
20101231,53400,1.5441,1.5442,1.5439,1.5439
20101231,53500,1.5438,1.544,1.5438,1.544
20101231,53600,1.544,1.544,1.5436,1.5437
20101231,53700,1.5438,1.5439,1.5438,1.5438
20101231,53800,1.5439,1.5439,1.5438,1.5438
20101231,53900,1.5437,1.5437,1.5432,1.5433
20101231,54000,1.5434,1.5437,1.5434,1.5436
20101231,54100,1.5436,1.5436,1.5434,1.5435
20101231,54200,1.5434,1.5435,1.5434,1.5435
20101231,54300,1.5435,1.5435,1.5434,1.5434
20101231,54400,1.5434,1.5434,1.5434,1.5434
20101231,54500,1.5433,1.5433,1.5432,1.5432
20101231,54600,1.5434,1.5435,1.5433,1.5434
20101231,54700,1.5435,1.5435,1.5433,1.5434
20101231,54800,1.5434,1.5435,1.5433,1.5435
20101231,54900,1.5436,1.5436,1.5435,1.5436
20101231,55000,1.5437,1.5437,1.5437,1.5437
20101231,55100,1.5437,1.5439,1.5436,1.5438
20101231,55200,1.5438,1.5438,1.5437,1.5437
20101231,55300,1.5437,1.5437,1.5436,1.5436
20101231,55400,1.5435,1.5438,1.5435,1.5436
20101231,55500,1.5437,1.5437,1.5435,1.5437
20101231,55600,1.5437,1.5437,1.5437,1.5437
20101231,55700,1.5437,1.5438,1.5437,1.5437
20101231,55800,1.5437,1.5437,1.5437,1.5437
20101231,55900,1.5437,1.5438,1.5437,1.5438
20101231,60000,1.5439,1.544,1.5439,1.544
20101231,60100,1.5439,1.5442,1.5439,1.5442
20101231,60200,1.5443,1.5443,1.5441,1.5441
20101231,60300,1.5441,1.5441,1.544,1.544
20101231,60400,1.544,1.5441,1.5439,1.544
20101231,60500,1.544,1.5441,1.5439,1.5439
20101231,60600,1.5439,1.5439,1.5437,1.5437
20101231,60700,1.5438,1.5441,1.5438,1.5441
20101231,60800,1.5441,1.5441,1.544,1.544
20101231,60900,1.544,1.544,1.544,1.544
20101231,61000,1.544,1.544,1.5438,1.544
20101231,61100,1.5441,1.5444,1.5441,1.5443
20101231,61200,1.5444,1.5444,1.544,1.5441
20101231,61300,1.5442,1.5449,1.5442,1.5447
20101231,61400,1.5446,1.5446,1.5445,1.5445
20101231,61500,1.5444,1.5445,1.5443,1.5443
20101231,61600,1.5443,1.5444,1.5442,1.5442
20101231,61700,1.5444,1.5444,1.5443,1.5443
20101231,61800,1.5443,1.5444,1.5442,1.5442
20101231,61900,1.5442,1.5442,1.5441,1.5442
20101231,62000,1.5444,1.5444,1.5442,1.5442
20101231,62100,1.5442,1.5444,1.5442,1.5443
20101231,62200,1.5444,1.5461,1.5444,1.5458
20101231,62300,1.5457,1.5459,1.5453,1.5459
20101231,62400,1.546,1.546,1.5453,1.5454
20101231,62500,1.5455,1.5456,1.5454,1.5455
20101231,62600,1.5454,1.5454,1.5453,1.5453
20101231,62700,1.5453,1.5454,1.5452,1.5454
20101231,62800,1.5454,1.5466,1.5454,1.5466
20101231,62900,1.5467,1.547,1.5461,1.5461
20101231,63000,1.546,1.5462,1.5454,1.546
20101231,63100,1.5459,1.5459,1.5457,1.5458
20101231,63200,1.5457,1.5457,1.545,1.545
20101231,63300,1.5449,1.5452,1.5448,1.5448
20101231,63400,1.5447,1.5454,1.5447,1.5454
20101231,63500,1.5455,1.546,1.5455,1.5458
20101231,63600,1.5458,1.5459,1.5457,1.5457
20101231,63700,1.5457,1.5461,1.5457,1.5461
20101231,63800,1.546,1.5463,1.546,1.5462
20101231,63900,1.5462,1.5462,1.5457,1.5457
20101231,64000,1.5458,1.5459,1.5458,1.5458
20101231,64100,1.5458,1.5458,1.5458,1.5458
20101231,64200,1.5458,1.5459,1.5456,1.5456
20101231,64300,1.5456,1.5456,1.5455,1.5456
20101231,64400,1.5456,1.5458,1.5456,1.5456
20101231,64500,1.5457,1.5458,1.5456,1.5458
20101231,64600,1.546,1.5466,1.546,1.5464
20101231,64700,1.5465,1.5465,1.5461,1.5463
20101231,64800,1.5464,1.5464,1.5462,1.5464
20101231,64900,1.5465,1.5469,1.5465,1.5469
20101231,65000,1.5468,1.5468,1.5464,1.5464
20101231,65100,1.5463,1.5463,1.5461,1.5462
20101231,65200,1.5463,1.5467,1.5463,1.5467
20101231,65300,1.5467,1.5476,1.5466,1.5476
20101231,65400,1.5475,1.5475,1.5473,1.5473
20101231,65500,1.5473,1.5474,1.5473,1.5474
20101231,65600,1.5474,1.5475,1.5474,1.5474
20101231,65700,1.5473,1.5474,1.5473,1.5474
20101231,65800,1.5474,1.5474,1.5473,1.5473
20101231,65900,1.5473,1.5474,1.5473,1.5474
20101231,70000,1.5474,1.5483,1.5474,1.5477
20101231,70100,1.5476,1.5481,1.5476,1.5479
20101231,70200,1.5478,1.5481,1.5478,1.5481
20101231,70300,1.5481,1.5483,1.5481,1.5483
20101231,70400,1.5482,1.5483,1.5481,1.5482
20101231,70500,1.5481,1.5481,1.5476,1.5476
20101231,70600,1.5475,1.5476,1.5475,1.5476
20101231,70700,1.5475,1.5476,1.5475,1.5476
20101231,70800,1.5477,1.5478,1.5477,1.5477
20101231,70900,1.5478,1.5478,1.5476,1.5476
20101231,71000,1.5476,1.5476,1.5473,1.5474
20101231,71100,1.5475,1.5478,1.5475,1.5475
20101231,71200,1.5476,1.5479,1.5476,1.5477
20101231,71300,1.5477,1.5477,1.5475,1.5476
20101231,71400,1.5476,1.5476,1.5475,1.5475
20101231,71500,1.5475,1.5476,1.5474,1.5474
20101231,71600,1.5473,1.5474,1.5472,1.5473
20101231,71700,1.5472,1.5473,1.5471,1.5471
20101231,71800,1.547,1.5472,1.5468,1.5472
20101231,71900,1.5472,1.5472,1.5472,1.5472
20101231,72000,1.5471,1.5474,1.5471,1.5474
20101231,72100,1.5474,1.5474,1.5473,1.5474
20101231,72200,1.5474,1.5474,1.5473,1.5473
20101231,72300,1.5472,1.5475,1.5472,1.5475
20101231,72400,1.5475,1.5484,1.5475,1.5484
20101231,72500,1.5486,1.549,1.5486,1.5489
20101231,72600,1.5488,1.5488,1.5483,1.5484
20101231,72700,1.5485,1.5485,1.548,1.5483
20101231,72800,1.5483,1.5484,1.5483,1.5483
20101231,72900,1.5484,1.5488,1.5484,1.5486
20101231,73000,1.5487,1.5487,1.5486,1.5487
20101231,73100,1.5487,1.5487,1.5485,1.5487
20101231,73200,1.5487,1.5488,1.5485,1.5486
20101231,73300,1.5485,1.5486,1.5484,1.5485
20101231,73400,1.5485,1.5485,1.5484,1.5484
20101231,73500,1.5483,1.5483,1.5481,1.5481
20101231,73600,1.5481,1.5484,1.5481,1.5483
20101231,73700,1.5482,1.5483,1.5482,1.5483
20101231,73800,1.5484,1.5484,1.5483,1.5483
20101231,73900,1.5482,1.5483,1.5482,1.5483
20101231,74000,1.5483,1.5484,1.5483,1.5484
20101231,74100,1.5484,1.5484,1.5482,1.5483
20101231,74200,1.5484,1.5485,1.5482,1.5483
20101231,74300,1.5484,1.5486,1.5484,1.5485
20101231,74400,1.5487,1.5491,1.5486,1.5486
20101231,74500,1.5485,1.5485,1.5483,1.5484
20101231,74600,1.5484,1.5486,1.5484,1.5486
20101231,74700,1.5486,1.5486,1.5483,1.5483
20101231,74800,1.5484,1.5486,1.5482,1.5485
20101231,74900,1.5486,1.5486,1.5485,1.5486
20101231,75000,1.5485,1.5488,1.5485,1.5487
20101231,75100,1.5488,1.5491,1.5488,1.5491
20101231,75200,1.5492,1.5496,1.5492,1.5495
20101231,75300,1.5496,1.5496,1.5495,1.5495
20101231,75400,1.5496,1.5496,1.5494,1.5496
20101231,75500,1.5496,1.5498,1.5495,1.5498
20101231,75600,1.5498,1.5499,1.5498,1.5499
20101231,75700,1.5499,1.5499,1.5498,1.5498
20101231,75800,1.5498,1.5498,1.5496,1.5496
20101231,75900,1.5495,1.5497,1.5494,1.5497
20101231,80000,1.5498,1.5504,1.5497,1.5504
20101231,80100,1.5505,1.5506,1.5502,1.5503
20101231,80200,1.5503,1.5504,1.5503,1.5503
20101231,80300,1.5502,1.5504,1.5502,1.5502
20101231,80400,1.5503,1.5504,1.55,1.55
20101231,80500,1.5499,1.5501,1.5499,1.5501
20101231,80600,1.5502,1.5502,1.5502,1.5502
20101231,80700,1.5501,1.5503,1.5498,1.5498
20101231,80800,1.5497,1.5497,1.5492,1.5492
20101231,80900,1.5492,1.5493,1.5492,1.5492
20101231,81000,1.5493,1.5493,1.5493,1.5493
20101231,81100,1.5493,1.5493,1.5488,1.5489
20101231,81200,1.5487,1.5488,1.5484,1.5488
20101231,81300,1.5488,1.5489,1.5487,1.5487
20101231,81400,1.5488,1.5489,1.5488,1.5488
20101231,81500,1.5488,1.5496,1.5487,1.5496
20101231,81600,1.5499,1.5503,1.5499,1.5503
20101231,81700,1.5502,1.5502,1.5495,1.5496
20101231,81800,1.5496,1.5496,1.5495,1.5495
20101231,81900,1.5495,1.5496,1.5494,1.5494
20101231,82000,1.5495,1.5497,1.5494,1.5496
20101231,82100,1.5495,1.5495,1.5494,1.5494
20101231,82200,1.5495,1.5495,1.5493,1.5493
20101231,82300,1.5493,1.5493,1.5493,1.5493
20101231,82400,1.5493,1.5493,1.5492,1.5492
20101231,82500,1.5491,1.5491,1.5484,1.5484
20101231,82600,1.5485,1.5485,1.5482,1.5484
20101231,82700,1.5484,1.5485,1.548,1.5485
20101231,82800,1.5486,1.5486,1.548,1.548
20101231,82900,1.5481,1.5482,1.5481,1.5482
20101231,83000,1.5483,1.5484,1.5482,1.5483
20101231,83100,1.5482,1.5483,1.5482,1.5482
20101231,83200,1.5481,1.5484,1.5481,1.5484
20101231,83300,1.5483,1.5484,1.5482,1.5482
20101231,83400,1.5482,1.5483,1.548,1.548
20101231,83500,1.5479,1.548,1.5474,1.5474
20101231,83600,1.5474,1.5474,1.547,1.547
20101231,83700,1.5471,1.5472,1.5468,1.5472
20101231,83800,1.5473,1.5474,1.5473,1.5474
20101231,83900,1.5475,1.5476,1.5473,1.5474
20101231,84000,1.5474,1.5474,1.5473,1.5474
20101231,84100,1.5474,1.5474,1.5473,1.5474
20101231,84200,1.5475,1.5476,1.5474,1.5474
20101231,84300,1.5473,1.5473,1.5471,1.5473
20101231,84400,1.5473,1.5482,1.5473,1.5479
20101231,84500,1.5479,1.5479,1.5475,1.5475
20101231,84600,1.5475,1.548,1.5475,1.548
20101231,84700,1.5481,1.5482,1.5478,1.5478
20101231,84800,1.5478,1.5478,1.5476,1.5476
20101231,84900,1.5477,1.5479,1.5477,1.5477
20101231,85000,1.5477,1.5479,1.5477,1.5479
20101231,85100,1.5478,1.5479,1.5477,1.5479
20101231,85200,1.5479,1.5479,1.5478,1.5479
20101231,85300,1.548,1.548,1.5478,1.5478
20101231,85400,1.5478,1.5478,1.5477,1.5477
20101231,85500,1.5478,1.548,1.5478,1.548
20101231,85600,1.5481,1.5482,1.5481,1.5482
20101231,85700,1.5482,1.5484,1.5481,1.5482
20101231,85800,1.5481,1.5481,1.5475,1.5475
20101231,85900,1.5475,1.5475,1.5474,1.5474
20101231,90000,1.5473,1.5473,1.547,1.5473
20101231,90100,1.5472,1.5478,1.547,1.5478
20101231,90200,1.5479,1.5479,1.5476,1.5477
20101231,90300,1.5478,1.5479,1.5473,1.5473
20101231,90400,1.5474,1.5478,1.5474,1.5476
20101231,90500,1.5477,1.5478,1.5474,1.5474
20101231,90600,1.5474,1.5474,1.5473,1.5473
20101231,90700,1.5473,1.5474,1.5473,1.5474
20101231,90800,1.5474,1.5474,1.5473,1.5474
20101231,90900,1.5474,1.5474,1.5472,1.5474
20101231,91000,1.5474,1.5475,1.5474,1.5474
20101231,91100,1.5473,1.5473,1.5468,1.5468
20101231,91200,1.5467,1.547,1.5467,1.547
20101231,91300,1.547,1.5473,1.547,1.5473
20101231,91400,1.5474,1.5474,1.5474,1.5474
20101231,91500,1.5474,1.5476,1.5474,1.5476
20101231,91600,1.5476,1.5477,1.5476,1.5477
20101231,91700,1.5476,1.5476,1.5475,1.5476
20101231,91800,1.5475,1.5475,1.5471,1.5471
20101231,91900,1.5472,1.5472,1.547,1.547
20101231,92000,1.547,1.547,1.5467,1.5467
20101231,92100,1.5467,1.5467,1.5467,1.5467
20101231,92200,1.5468,1.5468,1.5463,1.5463
20101231,92300,1.5462,1.5464,1.5461,1.5464
20101231,92400,1.5463,1.5466,1.5463,1.5464
20101231,92500,1.5463,1.5464,1.546,1.546
20101231,92600,1.546,1.546,1.5459,1.546
20101231,92700,1.5461,1.5468,1.5461,1.5468
20101231,92800,1.5468,1.5469,1.5467,1.5469
20101231,92900,1.5469,1.5469,1.5469,1.5469
20101231,93000,1.547,1.547,1.5469,1.547
20101231,93100,1.5469,1.5471,1.5468,1.547
20101231,93200,1.5469,1.5471,1.5469,1.5471
20101231,93300,1.5472,1.5472,1.547,1.5471
20101231,93400,1.547,1.5471,1.547,1.5471
20101231,93500,1.5472,1.5474,1.5472,1.5473
20101231,93600,1.5474,1.5477,1.5474,1.5477
20101231,93700,1.5478,1.5479,1.5478,1.5479
20101231,93800,1.548,1.548,1.5478,1.548
20101231,93900,1.548,1.5482,1.548,1.5482
20101231,94000,1.5483,1.5484,1.5478,1.5479
20101231,94100,1.548,1.548,1.5479,1.5479
20101231,94200,1.5479,1.548,1.5479,1.548
20101231,94300,1.5481,1.5482,1.5481,1.5482
20101231,94400,1.5482,1.5482,1.548,1.5482
20101231,94500,1.5482,1.5483,1.548,1.5483
20101231,94600,1.5484,1.5487,1.5484,1.5487
20101231,94700,1.5486,1.5489,1.5485,1.5489
20101231,94800,1.5488,1.5491,1.5488,1.549
20101231,94900,1.5491,1.5498,1.5491,1.5498
20101231,95000,1.5498,1.5498,1.5496,1.5497
20101231,95100,1.5497,1.5497,1.5496,1.5496
20101231,95200,1.5497,1.5498,1.5496,1.5497
20101231,95300,1.5498,1.5503,1.5497,1.5502
20101231,95400,1.5501,1.5501,1.5495,1.5495
20101231,95500,1.5495,1.5495,1.5495,1.5495
20101231,95600,1.5496,1.5496,1.5494,1.5495
20101231,95700,1.5495,1.5496,1.5495,1.5495
20101231,95800,1.5495,1.5495,1.5493,1.5495
20101231,95900,1.5494,1.5495,1.5494,1.5495
20101231,100000,1.5495,1.5496,1.5495,1.5495
20101231,100100,1.5494,1.5496,1.5494,1.5496
20101231,100200,1.5496,1.5496,1.5496,1.5496
20101231,100300,1.5496,1.5497,1.5496,1.5497
20101231,100400,1.5497,1.5497,1.5495,1.5495
20101231,100500,1.5495,1.5495,1.5494,1.5495
20101231,100600,1.5495,1.5496,1.5495,1.5496
20101231,100700,1.5496,1.5497,1.5496,1.5496
20101231,100800,1.5497,1.5497,1.5496,1.5496
20101231,100900,1.5496,1.5497,1.5495,1.5496
20101231,101000,1.5497,1.5497,1.5496,1.5496
20101231,101100,1.5497,1.5499,1.5497,1.5499
20101231,101200,1.5499,1.55,1.5496,1.5497
20101231,101300,1.5497,1.5497,1.5497,1.5497
20101231,101400,1.5496,1.5496,1.5495,1.5496
20101231,101500,1.5497,1.5497,1.5494,1.5494
20101231,101600,1.5495,1.5497,1.5495,1.5497
20101231,101700,1.5496,1.5496,1.5495,1.5495
20101231,101800,1.5496,1.5498,1.5495,1.5498
20101231,101900,1.5499,1.5503,1.5498,1.5503
20101231,102000,1.5502,1.5504,1.55,1.5504
20101231,102100,1.5505,1.5523,1.5505,1.5522
20101231,102200,1.5521,1.5521,1.5513,1.5514
20101231,102300,1.5513,1.5515,1.5513,1.5515
20101231,102400,1.5516,1.5519,1.5516,1.5518
20101231,102500,1.5517,1.5517,1.551,1.551
20101231,102600,1.5509,1.5511,1.5508,1.5508
20101231,102700,1.5509,1.5514,1.5509,1.5514
20101231,102800,1.5514,1.5517,1.5514,1.5517
20101231,102900,1.5516,1.5517,1.5516,1.5517
20101231,103000,1.5517,1.5517,1.5516,1.5516
20101231,103100,1.5517,1.5517,1.5516,1.5517
20101231,103200,1.5517,1.5518,1.5514,1.5518
20101231,103300,1.552,1.5525,1.552,1.5524
20101231,103400,1.5525,1.5527,1.5524,1.5525
20101231,103500,1.5524,1.5524,1.552,1.552
20101231,103600,1.552,1.552,1.5515,1.5519
20101231,103700,1.5518,1.5519,1.5516,1.5519
20101231,103800,1.5518,1.5519,1.5518,1.5518
20101231,103900,1.5517,1.5517,1.5515,1.5516
20101231,104000,1.5515,1.5516,1.5514,1.5515
20101231,104100,1.5516,1.5517,1.5515,1.5517
20101231,104200,1.5518,1.5518,1.5515,1.5515
20101231,104300,1.5514,1.5515,1.5514,1.5514
20101231,104400,1.5513,1.5513,1.5512,1.5512
20101231,104500,1.5513,1.5513,1.551,1.551
20101231,104600,1.5511,1.5511,1.5511,1.5511
20101231,104700,1.5511,1.5511,1.5509,1.551
20101231,104800,1.5511,1.5511,1.551,1.5511
20101231,104900,1.551,1.551,1.5502,1.5503
20101231,105000,1.5502,1.5504,1.5499,1.5504
20101231,105100,1.5503,1.5504,1.5501,1.5501
20101231,105200,1.5502,1.5503,1.5502,1.5502
20101231,105300,1.5503,1.5503,1.5498,1.5498
20101231,105400,1.5497,1.5497,1.5492,1.5493
20101231,105500,1.5492,1.5492,1.549,1.549
20101231,105600,1.5489,1.5494,1.5489,1.5493
20101231,105700,1.5491,1.5494,1.5491,1.5493
20101231,105800,1.5492,1.5492,1.549,1.549
20101231,105900,1.549,1.549,1.5486,1.5487
20101231,110000,1.5486,1.5486,1.5479,1.5485
20101231,110100,1.5484,1.5485,1.5482,1.5485
20101231,110200,1.5486,1.5487,1.5481,1.5481
20101231,110300,1.5482,1.5482,1.5482,1.5482
20101231,110400,1.5483,1.5483,1.5481,1.5482
20101231,110500,1.5481,1.5481,1.5481,1.5481
20101231,110600,1.5481,1.5481,1.5479,1.5481
20101231,110700,1.5481,1.5482,1.5481,1.5482
20101231,110800,1.5481,1.5484,1.5481,1.5482
20101231,110900,1.5482,1.5483,1.5481,1.5481
20101231,111000,1.548,1.5481,1.548,1.5481
20101231,111100,1.5481,1.5481,1.5481,1.5481
20101231,111200,1.5481,1.5481,1.5479,1.5479
20101231,111300,1.5479,1.5481,1.5479,1.548
20101231,111400,1.5479,1.548,1.5476,1.5476
20101231,111500,1.5477,1.5479,1.5477,1.5478
20101231,111600,1.5479,1.5481,1.5479,1.5481
20101231,111700,1.5481,1.5482,1.5481,1.5482
20101231,111800,1.5483,1.5485,1.5482,1.5484
20101231,111900,1.5483,1.5483,1.5482,1.5483
20101231,112000,1.5483,1.5483,1.5482,1.5483
20101231,112100,1.5482,1.5483,1.5482,1.5482
20101231,112200,1.5482,1.5483,1.5482,1.5483
20101231,112300,1.5483,1.5484,1.5483,1.5483
20101231,112400,1.5483,1.5487,1.5482,1.5482
20101231,112500,1.5482,1.5486,1.5482,1.5486
20101231,112600,1.5487,1.5489,1.5487,1.5488
20101231,112700,1.5488,1.5489,1.5488,1.5489
20101231,112800,1.5488,1.549,1.5488,1.549
20101231,112900,1.549,1.549,1.5486,1.5486
20101231,113000,1.5485,1.5487,1.5485,1.5487
20101231,113100,1.5487,1.5487,1.5485,1.5486
20101231,113200,1.5486,1.5491,1.5486,1.5491
20101231,113300,1.549,1.5492,1.549,1.5492
20101231,113400,1.5493,1.5494,1.5492,1.5492
20101231,113500,1.5491,1.5491,1.5489,1.549
20101231,113600,1.5491,1.5497,1.5489,1.5497
20101231,113700,1.5496,1.5496,1.5492,1.5495
20101231,113800,1.5496,1.5497,1.5496,1.5496
20101231,113900,1.5495,1.5501,1.5495,1.5499
20101231,114000,1.5498,1.5499,1.5497,1.5498
20101231,114100,1.5499,1.5503,1.5498,1.5503
20101231,114200,1.5502,1.5502,1.5501,1.5502
20101231,114300,1.5503,1.5506,1.5503,1.5506
20101231,114400,1.5505,1.5505,1.5503,1.5504
20101231,114500,1.5504,1.5504,1.5503,1.5504
20101231,114600,1.5504,1.5505,1.5504,1.5505
20101231,114700,1.5504,1.5505,1.5504,1.5505
20101231,114800,1.5504,1.5504,1.5502,1.5504
20101231,114900,1.5504,1.5504,1.5503,1.5504
20101231,115000,1.5504,1.5506,1.5503,1.5506
20101231,115100,1.5507,1.5511,1.5507,1.5511
20101231,115200,1.5512,1.5514,1.5512,1.5514
20101231,115300,1.5514,1.5515,1.5512,1.5515
20101231,115400,1.5516,1.5518,1.5515,1.5515
20101231,115500,1.5514,1.5514,1.5513,1.5513
20101231,115600,1.5512,1.5518,1.5512,1.5518
20101231,115700,1.5517,1.5522,1.5517,1.5522
20101231,115800,1.5523,1.5526,1.5522,1.5526
20101231,115900,1.5525,1.5525,1.5521,1.5521
20101231,120000,1.552,1.5528,1.5518,1.5525
20101231,120100,1.5526,1.5526,1.5519,1.5519
20101231,120200,1.552,1.5523,1.552,1.5523
20101231,120300,1.5522,1.5523,1.5522,1.5522
20101231,120400,1.5522,1.5523,1.5522,1.5522
20101231,120500,1.5521,1.5523,1.5521,1.5522
20101231,120600,1.5523,1.5524,1.5523,1.5523
20101231,120700,1.5522,1.5523,1.5521,1.5523
20101231,120800,1.5524,1.5524,1.5522,1.5524
20101231,120900,1.5523,1.5524,1.5523,1.5524
20101231,121000,1.5524,1.5524,1.5522,1.5523
20101231,121100,1.5523,1.5523,1.5522,1.5522
20101231,121200,1.5523,1.5524,1.5522,1.5522
20101231,121300,1.5521,1.5523,1.5521,1.5523
20101231,121400,1.5522,1.5524,1.5521,1.5524
20101231,121500,1.5523,1.5524,1.5523,1.5523
20101231,121600,1.5523,1.5524,1.5522,1.5522
20101231,121700,1.5523,1.5524,1.5522,1.5523
20101231,121800,1.5522,1.5522,1.5519,1.552
20101231,121900,1.5521,1.5523,1.5521,1.5521
20101231,122000,1.552,1.5524,1.552,1.5524
20101231,122100,1.5524,1.5525,1.5524,1.5525
20101231,122200,1.5524,1.5525,1.5524,1.5524
20101231,122300,1.5524,1.5524,1.5523,1.5524
20101231,122400,1.5524,1.5526,1.5524,1.5526
20101231,122500,1.5527,1.5527,1.5526,1.5527
20101231,122600,1.5527,1.5527,1.5527,1.5527
20101231,122700,1.5527,1.5527,1.5524,1.5524
20101231,122800,1.5523,1.5524,1.552,1.5523
20101231,122900,1.5523,1.5523,1.5522,1.5523
20101231,123000,1.5522,1.5523,1.5519,1.5519
20101231,123100,1.5519,1.5519,1.5515,1.5516
20101231,123200,1.5515,1.5522,1.5515,1.5522
20101231,123300,1.5522,1.5523,1.552,1.5523
20101231,123400,1.5522,1.5522,1.5517,1.552
20101231,123500,1.5521,1.5521,1.552,1.552
20101231,123600,1.5519,1.5523,1.5519,1.5523
20101231,123700,1.5524,1.5524,1.5522,1.5522
20101231,123800,1.5521,1.5523,1.552,1.5523
20101231,123900,1.5523,1.5527,1.5523,1.5526
20101231,124000,1.5527,1.5529,1.5527,1.5527
20101231,124100,1.5528,1.5529,1.5527,1.5527
20101231,124200,1.5528,1.553,1.5527,1.553
20101231,124300,1.5531,1.5532,1.5531,1.5531
20101231,124400,1.5532,1.5533,1.5531,1.5533
20101231,124500,1.5533,1.5536,1.5533,1.5535
20101231,124600,1.5536,1.5536,1.5536,1.5536
20101231,124700,1.5535,1.5541,1.5535,1.5541
20101231,124800,1.5542,1.5544,1.5539,1.554
20101231,124900,1.554,1.5541,1.5537,1.5537
20101231,125000,1.5538,1.5538,1.5528,1.5528
20101231,125100,1.5527,1.5527,1.5521,1.5521
20101231,125200,1.5521,1.5523,1.552,1.5523
20101231,125300,1.5523,1.5523,1.5523,1.5523
20101231,125400,1.5523,1.5523,1.5516,1.5517
20101231,125500,1.5518,1.5522,1.5518,1.5518
20101231,125600,1.5519,1.5522,1.5519,1.5521
20101231,125700,1.5521,1.5523,1.5521,1.5523
20101231,125800,1.5522,1.5522,1.5515,1.5516
20101231,125900,1.5516,1.5517,1.5516,1.5516
20101231,130000,1.5517,1.552,1.5517,1.552
20101231,130100,1.5521,1.5523,1.552,1.5521
20101231,130200,1.552,1.5524,1.5518,1.552
20101231,130300,1.5521,1.5523,1.552,1.5522
20101231,130400,1.5523,1.5524,1.5523,1.5524
20101231,130500,1.5523,1.5524,1.5522,1.5523
20101231,130600,1.5524,1.5524,1.5523,1.5523
20101231,130700,1.5523,1.5524,1.5523,1.5524
20101231,130800,1.5524,1.5525,1.5524,1.5524
20101231,130900,1.5525,1.5527,1.5525,1.5526
20101231,131000,1.5525,1.5525,1.5522,1.5524
20101231,131100,1.5525,1.5527,1.5525,1.5527
20101231,131200,1.5526,1.5529,1.5526,1.5528
20101231,131300,1.5528,1.5528,1.5528,1.5528
20101231,131400,1.5528,1.5529,1.5525,1.5525
20101231,131500,1.5525,1.5527,1.5522,1.5522
20101231,131600,1.5523,1.5523,1.5521,1.5522
20101231,131700,1.5521,1.5522,1.5521,1.5522
20101231,131800,1.5522,1.5523,1.5521,1.5523
20101231,131900,1.5524,1.5524,1.5523,1.5523
20101231,132000,1.5524,1.5528,1.5524,1.5528
20101231,132100,1.5527,1.5527,1.5525,1.5525
20101231,132200,1.5524,1.5528,1.5524,1.5527
20101231,132300,1.5528,1.5528,1.5526,1.5526
20101231,132400,1.5528,1.553,1.5528,1.5529
20101231,132500,1.5529,1.5529,1.5527,1.5528
20101231,132600,1.5529,1.5529,1.5527,1.5527
20101231,132700,1.5529,1.5531,1.5529,1.5531
20101231,132800,1.5532,1.5532,1.5532,1.5532
20101231,132900,1.5531,1.5531,1.5526,1.5526
20101231,133000,1.5525,1.5526,1.5525,1.5526
20101231,133100,1.5526,1.5526,1.5524,1.5524
20101231,133200,1.5523,1.5524,1.5521,1.5521
20101231,133300,1.552,1.5522,1.5519,1.5522
20101231,133400,1.5521,1.5522,1.552,1.552
20101231,133500,1.5519,1.552,1.5519,1.552
20101231,133600,1.552,1.552,1.5519,1.5519
20101231,133700,1.552,1.552,1.5516,1.5517
20101231,133800,1.5518,1.5519,1.5518,1.5519
20101231,133900,1.552,1.5524,1.552,1.5523
20101231,134000,1.5524,1.5524,1.5521,1.5522
20101231,134100,1.5521,1.5523,1.5521,1.5523
20101231,134200,1.5523,1.5524,1.5523,1.5524
20101231,134300,1.5524,1.5524,1.5523,1.5524
20101231,134400,1.5524,1.5524,1.5523,1.5523
20101231,134500,1.5522,1.5522,1.5521,1.5521
20101231,134600,1.5521,1.5521,1.5519,1.5519
20101231,134700,1.552,1.5522,1.5519,1.552
20101231,134800,1.5521,1.5521,1.5519,1.5519
20101231,134900,1.5519,1.5519,1.5515,1.5515
20101231,135000,1.5516,1.5518,1.5514,1.5514
20101231,135100,1.5514,1.5518,1.5514,1.5518
20101231,135200,1.5519,1.5525,1.5519,1.5525
20101231,135300,1.5526,1.5528,1.5525,1.5525
20101231,135400,1.5524,1.5524,1.5523,1.5523
20101231,135500,1.5521,1.5523,1.5521,1.5523
20101231,135600,1.5522,1.5523,1.5522,1.5522
20101231,135700,1.5521,1.5521,1.5519,1.5519
20101231,135800,1.5518,1.552,1.5518,1.552
20101231,135900,1.552,1.552,1.5518,1.5519
20101231,140000,1.5518,1.5519,1.5518,1.5519
20101231,140100,1.5519,1.5519,1.5518,1.5519
20101231,140200,1.5518,1.5521,1.5518,1.5521
20101231,140300,1.552,1.5521,1.552,1.552
20101231,140400,1.552,1.5521,1.552,1.5521
20101231,140500,1.5522,1.5522,1.552,1.5521
20101231,140600,1.552,1.5523,1.552,1.5523
20101231,140700,1.5523,1.5525,1.5523,1.5525
20101231,140800,1.5525,1.5525,1.5525,1.5525
20101231,140900,1.5525,1.5525,1.5522,1.5524
20101231,141000,1.5524,1.5524,1.5524,1.5524
20101231,141100,1.5525,1.5525,1.5524,1.5524
20101231,141200,1.5525,1.5528,1.5525,1.5528
20101231,141300,1.5527,1.5527,1.5525,1.5525
20101231,141400,1.5524,1.5528,1.5524,1.5528
20101231,141500,1.5529,1.5532,1.5528,1.5532
20101231,141600,1.5531,1.5533,1.553,1.5532
20101231,141700,1.5531,1.5531,1.553,1.553
20101231,141800,1.553,1.553,1.5529,1.5529
20101231,141900,1.553,1.553,1.5529,1.5529
20101231,142000,1.5529,1.553,1.5528,1.5528
20101231,142100,1.5529,1.5529,1.5526,1.5527
20101231,142200,1.5528,1.5529,1.5528,1.5529
20101231,142300,1.5529,1.5531,1.5527,1.5531
20101231,142400,1.5532,1.5545,1.5531,1.5545
20101231,142500,1.5544,1.5545,1.5541,1.5541
20101231,142600,1.554,1.5541,1.5539,1.5539
20101231,142700,1.5538,1.5542,1.5538,1.5541
20101231,142800,1.554,1.554,1.5539,1.5539
20101231,142900,1.5541,1.5541,1.554,1.5541
20101231,143000,1.5541,1.5543,1.554,1.5543
20101231,143100,1.5544,1.5549,1.5544,1.5549
20101231,143200,1.555,1.5555,1.555,1.5553
20101231,143300,1.5554,1.5559,1.5554,1.5558
20101231,143400,1.5559,1.5575,1.5559,1.5572
20101231,143500,1.5571,1.5578,1.5569,1.557
20101231,143600,1.557,1.5572,1.557,1.557
20101231,143700,1.5571,1.5572,1.5571,1.5572
20101231,143800,1.5573,1.5578,1.5573,1.5578
20101231,143900,1.5578,1.5582,1.5578,1.5581
20101231,144000,1.558,1.5581,1.5577,1.5577
20101231,144100,1.5576,1.5579,1.5576,1.5579
20101231,144200,1.5579,1.5584,1.5579,1.5583
20101231,144300,1.5583,1.5583,1.558,1.5581
20101231,144400,1.5582,1.5582,1.558,1.558
20101231,144500,1.5581,1.5581,1.5579,1.558
20101231,144600,1.5579,1.5579,1.5577,1.5578
20101231,144700,1.5579,1.5581,1.5579,1.5581
20101231,144800,1.5582,1.5583,1.5576,1.5576
20101231,144900,1.5575,1.5576,1.5575,1.5576
20101231,145000,1.5576,1.5576,1.5574,1.5576
20101231,145100,1.5578,1.5578,1.5576,1.5576
20101231,145200,1.5576,1.5577,1.5575,1.5576
20101231,145300,1.5575,1.5576,1.5574,1.5576
20101231,145400,1.5576,1.5581,1.5576,1.5581
20101231,145500,1.5582,1.5584,1.5581,1.5581
20101231,145600,1.5582,1.5582,1.5581,1.5582
20101231,145700,1.5581,1.5582,1.5581,1.5581
20101231,145800,1.5581,1.5582,1.558,1.558
20101231,145900,1.5579,1.558,1.5578,1.558
20101231,150000,1.5581,1.5581,1.5574,1.5574
20101231,150100,1.5573,1.5577,1.557,1.5577
20101231,150200,1.5577,1.5583,1.5577,1.5583
20101231,150300,1.5582,1.5583,1.5582,1.5582
20101231,150400,1.5582,1.5582,1.5582,1.5582
20101231,150500,1.5581,1.5582,1.5581,1.5582
20101231,150600,1.5582,1.5584,1.5582,1.5584
20101231,150700,1.5584,1.5584,1.5583,1.5584
20101231,150800,1.5585,1.5594,1.5585,1.5594
20101231,150900,1.5595,1.5601,1.5595,1.56
20101231,151000,1.5599,1.5599,1.5596,1.5596
20101231,151100,1.5595,1.5599,1.5594,1.5599
20101231,151200,1.56,1.5602,1.5596,1.5597
20101231,151300,1.5598,1.5599,1.5598,1.5598
20101231,151400,1.5597,1.5597,1.5595,1.5596
20101231,151500,1.5595,1.5595,1.5594,1.5594
20101231,151600,1.5594,1.5594,1.5592,1.5592
20101231,151700,1.5592,1.5592,1.5591,1.5591
20101231,151800,1.5591,1.5592,1.5589,1.5589
20101231,151900,1.559,1.559,1.5586,1.5587
20101231,152000,1.5588,1.559,1.5588,1.559
20101231,152100,1.5591,1.5591,1.5589,1.5589
20101231,152200,1.5588,1.559,1.5588,1.559
20101231,152300,1.5589,1.559,1.5589,1.5589
20101231,152400,1.5588,1.5592,1.5588,1.5592
20101231,152500,1.5593,1.5595,1.5591,1.5592
20101231,152600,1.5592,1.5596,1.5591,1.5594
20101231,152700,1.5595,1.56,1.5595,1.56
20101231,152800,1.5599,1.5604,1.5599,1.5604
20101231,152900,1.5603,1.5605,1.5603,1.5605
20101231,153000,1.5605,1.5605,1.5603,1.5603
20101231,153100,1.5603,1.5603,1.5603,1.5603
20101231,153200,1.5603,1.5603,1.5602,1.5602
20101231,153300,1.5602,1.5602,1.56,1.5601
20101231,153400,1.56,1.5602,1.56,1.5602
20101231,153500,1.5603,1.5611,1.5603,1.5611
20101231,153600,1.5612,1.5613,1.5612,1.5612
20101231,153700,1.5613,1.5616,1.5613,1.5616
20101231,153800,1.5617,1.5622,1.5616,1.5622
20101231,153900,1.5621,1.5621,1.562,1.5621
20101231,154000,1.5622,1.5627,1.5622,1.5627
20101231,154100,1.5627,1.5627,1.5623,1.5625
20101231,154200,1.5625,1.5625,1.5624,1.5625
20101231,154300,1.5626,1.563,1.5626,1.563
20101231,154400,1.5631,1.5634,1.563,1.5634
20101231,154500,1.5633,1.5634,1.5632,1.5634
20101231,154600,1.5634,1.5634,1.5626,1.5626
20101231,154700,1.5625,1.5625,1.5622,1.5623
20101231,154800,1.5623,1.5624,1.5623,1.5624
20101231,154900,1.5623,1.5627,1.5623,1.5627
20101231,155000,1.5628,1.5629,1.5627,1.5628
20101231,155100,1.5628,1.5629,1.5624,1.5624
20101231,155200,1.5625,1.5626,1.5623,1.5625
20101231,155300,1.5626,1.5631,1.5625,1.5631
20101231,155400,1.5632,1.5644,1.5632,1.5644
20101231,155500,1.5645,1.5649,1.5645,1.5649
20101231,155600,1.565,1.5652,1.5646,1.5646
20101231,155700,1.5647,1.5653,1.5647,1.5652
20101231,155800,1.5653,1.5653,1.5646,1.5647
20101231,155900,1.5648,1.5653,1.5648,1.5652
20101231,160000,1.5651,1.5662,1.5648,1.5657
20101231,160100,1.5655,1.5655,1.5638,1.5641
20101231,160200,1.5642,1.5647,1.5642,1.5643
20101231,160300,1.5644,1.5647,1.5644,1.5647
20101231,160400,1.5646,1.5647,1.5645,1.5647
20101231,160500,1.5646,1.5646,1.5644,1.5645
20101231,160600,1.5646,1.5648,1.5644,1.5644
20101231,160700,1.5643,1.5643,1.5631,1.5633
20101231,160800,1.5634,1.5635,1.5633,1.5634
20101231,160900,1.5635,1.5635,1.5634,1.5634
20101231,161000,1.5634,1.5634,1.5628,1.5628
20101231,161100,1.5627,1.5627,1.562,1.562
20101231,161200,1.5619,1.5619,1.5616,1.5616
20101231,161300,1.5616,1.562,1.5616,1.5619
20101231,161400,1.562,1.562,1.5616,1.5617
20101231,161500,1.5618,1.5618,1.5602,1.5604
20101231,161600,1.5604,1.5605,1.5604,1.5605
20101231,161700,1.5604,1.5605,1.5604,1.5605
20101231,161800,1.5605,1.5606,1.5604,1.5606
20101231,161900,1.5605,1.5606,1.5605,1.5606
20101231,162000,1.5607,1.5609,1.5607,1.5608
20101231,162100,1.5608,1.5609,1.5608,1.5608
20101231,162200,1.5607,1.5615,1.5607,1.5614
20101231,162300,1.5613,1.5617,1.5611,1.5616
20101231,162400,1.5617,1.5617,1.5611,1.5611
20101231,162500,1.5611,1.5616,1.561,1.5615
20101231,162600,1.5614,1.5614,1.5603,1.5604
20101231,162700,1.5605,1.5608,1.5605,1.5607
20101231,162800,1.5608,1.5609,1.5605,1.5605
20101231,162900,1.5605,1.5607,1.5604,1.5604
20101231,163000,1.5605,1.5612,1.5605,1.5612
20101231,163100,1.5613,1.5616,1.5613,1.5613
20101231,163200,1.5613,1.5614,1.5609,1.5609
20101231,163300,1.5608,1.5608,1.5607,1.5607
20101231,163400,1.5607,1.5608,1.5607,1.5607
20101231,163500,1.5608,1.561,1.5608,1.561
20101231,163600,1.561,1.5615,1.561,1.5614
20101231,163700,1.5613,1.5615,1.5613,1.5613
20101231,163800,1.5613,1.5613,1.5611,1.5612
20101231,163900,1.5612,1.5614,1.5611,1.5613
20101231,164000,1.5614,1.5617,1.5614,1.5617
20101231,164100,1.5616,1.5617,1.5615,1.5616
20101231,164200,1.5616,1.5616,1.5616,1.5616
20101231,164300,1.5617,1.562,1.5617,1.5618
20101231,164400,1.5618,1.5619,1.5618,1.5619
20101231,164500,1.5619,1.5619,1.5615,1.5615
20101231,164600,1.5614,1.5615,1.5614,1.5614
20101231,164700,1.5614,1.5614,1.5614,1.5614
20101231,164800,1.5614,1.5614,1.5612,1.5612
20101231,164900,1.5611,1.5613,1.5611,1.5613
20101231,165000,1.5612,1.5612,1.5607,1.5607
20101231,165100,1.5608,1.5612,1.5608,1.5612
20101231,165200,1.5612,1.5612,1.5611,1.5611
20101231,165300,1.561,1.5612,1.561,1.5611
20101231,165400,1.561,1.5614,1.561,1.5614
20101231,165500,1.5615,1.5616,1.5615,1.5616
20101231,165600,1.5617,1.5617,1.5616,1.5616
20101231,165700,1.5616,1.5616,1.5614,1.5614
20101231,165800,1.5613,1.5613,1.5609,1.5609
20101231,165900,1.561,1.561,1.5605,1.5606
20101231,170000,1.5605,1.5605,1.5595,1.5595
20101231,170100,1.5594,1.5594,1.5593,1.5593
20101231,170200,1.5594,1.5594,1.5593,1.5594
20101231,170300,1.5594,1.5595,1.5594,1.5595
20101231,170400,1.5595,1.5599,1.5595,1.5597
20101231,170500,1.5597,1.5597,1.5594,1.5594
20101231,170600,1.5593,1.5594,1.5592,1.5594
20101231,170700,1.5595,1.5595,1.5591,1.5594
20101231,170800,1.5595,1.5599,1.5594,1.5599
20101231,170900,1.5601,1.5602,1.5601,1.5602
20101231,171000,1.5603,1.5605,1.5603,1.5605
20101231,171100,1.5606,1.5606,1.5605,1.5605
20101231,171200,1.5604,1.5604,1.5599,1.5601
20101231,171300,1.5603,1.5606,1.5602,1.5606
20101231,171400,1.5605,1.5608,1.5605,1.5608
20101231,171500,1.561,1.5613,1.561,1.5613
20101231,171600,1.5612,1.5613,1.5611,1.5611
20101231,171700,1.5611,1.5611,1.5611,1.5611
20101231,171800,1.5612,1.5612,1.561,1.561
20101231,171900,1.5609,1.5609,1.5607,1.5607
20101231,172000,1.5608,1.5608,1.5607,1.5607
20101231,172100,1.5607,1.5608,1.5607,1.5607
20101231,172200,1.5607,1.5608,1.5607,1.5608
20101231,172300,1.5608,1.5608,1.5606,1.5606
20101231,172400,1.5607,1.5607,1.5605,1.5607
20101231,172500,1.5608,1.5611,1.5607,1.5611
20101231,172600,1.5612,1.5612,1.561,1.561
20101231,172700,1.5611,1.5615,1.5611,1.5612
20101231,172800,1.5611,1.5611,1.5611,1.5611
20101231,172900,1.5612,1.5612,1.5611,1.5612
20101231,173000,1.5611,1.5617,1.5611,1.5617
20101231,173100,1.5616,1.5617,1.5616,1.5617
20101231,173200,1.5616,1.5622,1.5615,1.5619
20101231,173300,1.5618,1.5618,1.5616,1.5617
20101231,173400,1.5616,1.5617,1.5616,1.5616
20101231,173500,1.5617,1.5617,1.5616,1.5616
20101231,173600,1.5615,1.5616,1.5614,1.5614
20101231,173700,1.5615,1.5616,1.5614,1.5615
20101231,173800,1.5614,1.5615,1.5613,1.5613
20101231,173900,1.5613,1.5613,1.5613,1.5613
20101231,174000,1.5614,1.5614,1.5611,1.5612
20101231,174100,1.5613,1.5615,1.5612,1.5614
20101231,174200,1.5614,1.5615,1.5614,1.5614
20101231,174300,1.5614,1.5615,1.5614,1.5614
20101231,174400,1.5614,1.5615,1.5613,1.5613
20101231,174500,1.5612,1.5612,1.5606,1.5607
20101231,174600,1.5606,1.5608,1.5606,1.5608
20101231,174700,1.5609,1.5609,1.5607,1.5608
20101231,174800,1.5608,1.5608,1.5608,1.5608
20101231,174900,1.5608,1.5609,1.5608,1.5609
20101231,175000,1.5609,1.5609,1.5608,1.5608
20101231,175100,1.5608,1.5608,1.5607,1.5608
20101231,175200,1.5607,1.5607,1.5604,1.5604
20101231,175300,1.5605,1.5605,1.5604,1.5605
20101231,175400,1.5605,1.5605,1.5604,1.5604
20101231,175500,1.5604,1.5604,1.5599,1.56
20101231,175600,1.5599,1.5599,1.5595,1.5596
20101231,175700,1.5595,1.5595,1.5594,1.5594
20101231,175800,1.5594,1.5595,1.5593,1.5593
20101231,175900,1.5592,1.5592,1.559,1.559
20101231,180000,1.5591,1.5591,1.5588,1.5588
20101231,180100,1.5587,1.5587,1.5583,1.5584
20101231,180200,1.5583,1.5585,1.5583,1.5584
20101231,180300,1.5583,1.5583,1.5583,1.5583
20101231,180400,1.5582,1.5582,1.5575,1.5576
20101231,180500,1.5577,1.5584,1.5577,1.5583
20101231,180600,1.5584,1.5588,1.5584,1.5586
20101231,180700,1.5586,1.5586,1.5585,1.5585
20101231,180800,1.5584,1.5585,1.5584,1.5585
20101231,180900,1.5585,1.5588,1.5585,1.5586
20101231,181000,1.5587,1.5588,1.5586,1.5588
20101231,181100,1.5589,1.5589,1.5588,1.5588
20101231,181200,1.5588,1.5588,1.5581,1.5584
20101231,181300,1.5583,1.5583,1.5581,1.5581
20101231,181400,1.5582,1.5584,1.5582,1.5584
20101231,181500,1.5584,1.5584,1.5582,1.5582
20101231,181600,1.5581,1.5581,1.5576,1.5576
20101231,181700,1.5577,1.558,1.5577,1.5579
20101231,181800,1.5577,1.5583,1.5577,1.5577
20101231,181900,1.5576,1.5576,1.5575,1.5575
20101231,182000,1.5574,1.5574,1.5572,1.5572
20101231,182100,1.5571,1.5571,1.557,1.557
20101231,182200,1.5571,1.5572,1.5571,1.5572
20101231,182300,1.5571,1.5571,1.5571,1.5571
20101231,182400,1.5571,1.5571,1.5571,1.5571
20101231,182500,1.5572,1.5572,1.5571,1.5572
20101231,182600,1.5573,1.5574,1.5573,1.5574
20101231,182700,1.5573,1.5574,1.5573,1.5574
20101231,182800,1.5575,1.5575,1.5574,1.5574
20101231,182900,1.5574,1.5574,1.5574,1.5574
20101231,183000,1.5575,1.5576,1.5575,1.5575
20101231,183100,1.5575,1.5577,1.5575,1.5577
20101231,183200,1.5576,1.5578,1.5576,1.5578
20101231,183300,1.5579,1.5579,1.5579,1.5579
20101231,183400,1.5578,1.5578,1.5575,1.5575
20101231,183500,1.5574,1.5576,1.5574,1.5575
20101231,183600,1.5574,1.5574,1.5574,1.5574
20101231,183700,1.5574,1.5574,1.5574,1.5574
20101231,183800,1.5574,1.5575,1.5574,1.5575
20101231,183900,1.5576,1.5576,1.5575,1.5575
20101231,184000,1.5575,1.5575,1.5575,1.5575
20101231,184100,1.5575,1.5575,1.5575,1.5575
20101231,184200,1.5575,1.5575,1.5575,1.5575
20101231,184300,1.5575,1.5575,1.5575,1.5575
20101231,184400,1.5575,1.5576,1.5575,1.5576
20101231,184500,1.5576,1.5576,1.5573,1.5573
20101231,184600,1.5572,1.5573,1.5572,1.5572
20101231,184700,1.5572,1.5572,1.5571,1.5572
20101231,184800,1.5573,1.5573,1.557,1.557
20101231,184900,1.5569,1.5569,1.5568,1.5568
20101231,185000,1.5569,1.5569,1.5568,1.5569
20101231,185100,1.5569,1.557,1.5569,1.557
20101231,185200,1.557,1.5571,1.5569,1.5571
20101231,185300,1.5571,1.5571,1.5571,1.5571
20101231,185400,1.557,1.557,1.5569,1.5569
20101231,185500,1.5569,1.5569,1.5565,1.5565
20101231,185600,1.5566,1.5566,1.5565,1.5565
20101231,185700,1.5565,1.5566,1.5565,1.5566
20101231,185800,1.5566,1.5566,1.5565,1.5566
20101231,185900,1.5566,1.5566,1.5565,1.5566
20101231,190000,1.5567,1.5567,1.5566,1.5566
20101231,190100,1.5566,1.5566,1.5566,1.5566
20101231,190200,1.5567,1.5567,1.5566,1.5566
20101231,190300,1.5566,1.5566,1.5566,1.5566
20101231,190400,1.5565,1.5565,1.5564,1.5565
20101231,190500,1.5565,1.5566,1.5565,1.5566
20101231,190600,1.5565,1.5566,1.5565,1.5565
20101231,190700,1.5565,1.5565,1.5564,1.5564
20101231,190800,1.5564,1.5565,1.5563,1.5563
20101231,190900,1.5562,1.5562,1.5557,1.556
20101231,191000,1.5558,1.5558,1.5556,1.5557
20101231,191100,1.5558,1.5558,1.5558,1.5558
20101231,191200,1.5558,1.5572,1.5557,1.5572
20101231,191300,1.5571,1.5571,1.5571,1.5571
20101231,191400,1.5571,1.5571,1.557,1.557
20101231,191500,1.557,1.5571,1.5569,1.5571
20101231,191600,1.5571,1.5571,1.5571,1.5571
20101231,191700,1.5571,1.5571,1.5571,1.5571
20101231,191800,1.5571,1.5571,1.557,1.5571
20101231,191900,1.5571,1.5571,1.557,1.5571
20101231,192000,1.5571,1.5571,1.557,1.557
20101231,192100,1.5569,1.557,1.5569,1.557
20101231,192200,1.557,1.5571,1.557,1.557
20101231,192300,1.557,1.557,1.557,1.557
20101231,192400,1.557,1.5571,1.557,1.5571
20101231,192500,1.5571,1.5571,1.5569,1.5569
20101231,192600,1.557,1.557,1.5569,1.5569
20101231,192700,1.5569,1.5569,1.5569,1.5569
20101231,192800,1.5569,1.5569,1.5566,1.5568
20101231,192900,1.5567,1.5567,1.5565,1.5565
20101231,193000,1.5564,1.5567,1.5564,1.5565
20101231,193100,1.5565,1.5565,1.5565,1.5565
20101231,193200,1.5565,1.5566,1.5565,1.5566
20101231,193300,1.5565,1.5567,1.5565,1.5567
20101231,193400,1.5567,1.5567,1.5566,1.5566
20101231,193500,1.5567,1.5567,1.5565,1.5565
20101231,193600,1.5564,1.5566,1.5564,1.5565
20101231,193700,1.5565,1.5565,1.5565,1.5565
20101231,193800,1.5565,1.5565,1.5565,1.5565
20101231,193900,1.5566,1.5566,1.5566,1.5566
20101231,194000,1.5566,1.5566,1.5565,1.5565
20101231,194100,1.5565,1.5565,1.5565,1.5565
20101231,194200,1.5565,1.5566,1.5565,1.5566
20101231,194300,1.5566,1.5566,1.5566,1.5566
20101231,194400,1.5566,1.5567,1.5566,1.5567
20101231,194500,1.5567,1.5567,1.5567,1.5567
20101231,194600,1.5567,1.5567,1.5566,1.5566
20101231,194700,1.5566,1.5569,1.5566,1.5568
20101231,194800,1.5569,1.5572,1.5569,1.5572
20101231,194900,1.5571,1.5572,1.5571,1.5572
20101231,195000,1.5573,1.5573,1.5573,1.5573
20101231,195100,1.5573,1.5573,1.5573,1.5573
20101231,195200,1.5573,1.5574,1.5573,1.5574
20101231,195300,1.5575,1.5583,1.5575,1.5583
20101231,195400,1.5583,1.5583,1.5582,1.5582
20101231,195500,1.5582,1.5585,1.5582,1.5585
20101231,195600,1.5586,1.5597,1.5586,1.5597
20101231,195700,1.5598,1.5619,1.5578,1.5584
20101231,195800,1.5585,1.5588,1.5584,1.5588
20101231,195900,1.5589,1.5589,1.5586,1.5586
20101231,200000,1.5587,1.559,1.5587,1.5589
20101231,200100,1.559,1.5594,1.559,1.5593
20101231,200200,1.5593,1.5595,1.5593,1.5595
20101231,200300,1.5594,1.5594,1.5592,1.5593
20101231,200400,1.5594,1.5594,1.5594,1.5594
20101231,200500,1.5593,1.5593,1.5593,1.5593
20101231,200600,1.5593,1.5594,1.559,1.559
20101231,200700,1.5594,1.5597,1.5594,1.5596
20101231,200800,1.5597,1.5597,1.5595,1.5595
20101231,200900,1.5597,1.5597,1.5596,1.5596
20101231,201000,1.5597,1.5597,1.5595,1.5595
20101231,201100,1.5596,1.5597,1.5596,1.5596
20101231,201200,1.5595,1.5595,1.5595,1.5595
20101231,201300,1.5596,1.5596,1.5595,1.5595
20101231,201400,1.5593,1.5593,1.5593,1.5593
20101231,201500,1.5593,1.5596,1.5593,1.5596
20101231,201600,1.5596,1.5596,1.5596,1.5596
20101231,201700,1.5596,1.5597,1.5596,1.5597
20101231,201800,1.5597,1.5599,1.5597,1.5599
20101231,201900,1.5599,1.5599,1.5599,1.5599
20101231,202000,1.5599,1.5599,1.5599,1.5599
20101231,202100,1.5603,1.5603,1.5601,1.5601
20101231,202200,1.5601,1.5604,1.5601,1.5604
20101231,202300,1.5606,1.5608,1.5603,1.5603
20101231,202400,1.5603,1.5603,1.5603,1.5603
20101231,202500,1.5603,1.5603,1.5603,1.5603
20101231,202600,1.5605,1.5605,1.5604,1.5604
20101231,202700,1.5604,1.5604,1.5604,1.5604
20101231,202800,1.5604,1.5604,1.5603,1.5603
20101231,202900,1.5603,1.5604,1.5603,1.5604
20101231,203000,1.5604,1.5604,1.5602,1.5602
20101231,203100,1.5603,1.5603,1.5601,1.5603
20101231,203200,1.5605,1.5605,1.5603,1.5603
20101231,203300,1.5604,1.5605,1.5604,1.5605
20101231,203400,1.5605,1.5607,1.5605,1.5607
20101231,203500,1.5607,1.5608,1.5605,1.5607
20101231,203600,1.5607,1.5608,1.5607,1.5608
20101231,203700,1.5608,1.5608,1.5607,1.5607
20101231,203800,1.5607,1.5607,1.5607,1.5607
20101231,203900,1.5606,1.5606,1.5602,1.5603
20101231,204000,1.5603,1.5603,1.5603,1.5603
20101231,204100,1.5603,1.5604,1.5603,1.5604
20101231,204200,1.5604,1.5605,1.5603,1.5603
20101231,204300,1.5604,1.5604,1.5602,1.5602
20101231,204400,1.5601,1.5601,1.5601,1.5601
20101231,204500,1.5601,1.5601,1.5601,1.5601
20101231,204600,1.5601,1.5601,1.5601,1.5601
20101231,204700,1.5601,1.5601,1.5599,1.5599
20101231,204800,1.5599,1.5599,1.5599,1.5599
20101231,204900,1.5599,1.5599,1.5599,1.5599
20101231,205000,1.5599,1.5599,1.5596,1.5596
20101231,205100,1.5595,1.5596,1.5595,1.5596
20101231,205200,1.5597,1.5597,1.5597,1.5597
20101231,205300,1.5597,1.5598,1.5597,1.5598
20101231,205400,1.5599,1.5599,1.5599,1.5599
20101231,205500,1.5599,1.5599,1.5598,1.5599
20101231,205600,1.5599,1.5599,1.5593,1.5593
20101231,205700,1.5592,1.5592,1.5591,1.5591
20101231,205800,1.5591,1.5591,1.5591,1.5591
20101231,205900,1.5591,1.5592,1.5591,1.5592
